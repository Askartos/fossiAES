magic
tech sky130A
magscale 1 2
timestamp 1653875649
<< obsli1 >>
rect 1104 2159 98808 97393
<< obsm1 >>
rect 14 2128 99898 97424
<< metal2 >>
rect 2594 99200 2650 100000
rect 8390 99200 8446 100000
rect 14830 99200 14886 100000
rect 20626 99200 20682 100000
rect 27066 99200 27122 100000
rect 32862 99200 32918 100000
rect 39302 99200 39358 100000
rect 45098 99200 45154 100000
rect 51538 99200 51594 100000
rect 57334 99200 57390 100000
rect 63774 99200 63830 100000
rect 69570 99200 69626 100000
rect 76010 99200 76066 100000
rect 81806 99200 81862 100000
rect 88246 99200 88302 100000
rect 94042 99200 94098 100000
rect 99838 99200 99894 100000
rect 18 0 74 800
rect 5814 0 5870 800
rect 11610 0 11666 800
rect 18050 0 18106 800
rect 23846 0 23902 800
rect 30286 0 30342 800
rect 36082 0 36138 800
rect 42522 0 42578 800
rect 48318 0 48374 800
rect 54758 0 54814 800
rect 60554 0 60610 800
rect 66994 0 67050 800
rect 72790 0 72846 800
rect 79230 0 79286 800
rect 85026 0 85082 800
rect 91466 0 91522 800
rect 97262 0 97318 800
<< obsm2 >>
rect 20 99144 2538 99362
rect 2706 99144 8334 99362
rect 8502 99144 14774 99362
rect 14942 99144 20570 99362
rect 20738 99144 27010 99362
rect 27178 99144 32806 99362
rect 32974 99144 39246 99362
rect 39414 99144 45042 99362
rect 45210 99144 51482 99362
rect 51650 99144 57278 99362
rect 57446 99144 63718 99362
rect 63886 99144 69514 99362
rect 69682 99144 75954 99362
rect 76122 99144 81750 99362
rect 81918 99144 88190 99362
rect 88358 99144 93986 99362
rect 94154 99144 99782 99362
rect 20 856 99892 99144
rect 130 800 5758 856
rect 5926 800 11554 856
rect 11722 800 17994 856
rect 18162 800 23790 856
rect 23958 800 30230 856
rect 30398 800 36026 856
rect 36194 800 42466 856
rect 42634 800 48262 856
rect 48430 800 54702 856
rect 54870 800 60498 856
rect 60666 800 66938 856
rect 67106 800 72734 856
rect 72902 800 79174 856
rect 79342 800 84970 856
rect 85138 800 91410 856
rect 91578 800 97206 856
rect 97374 800 99892 856
<< metal3 >>
rect 0 96568 800 96688
rect 99200 93168 100000 93288
rect 0 89768 800 89888
rect 99200 87048 100000 87168
rect 0 83648 800 83768
rect 99200 80248 100000 80368
rect 0 76848 800 76968
rect 99200 74128 100000 74248
rect 0 70728 800 70848
rect 99200 67328 100000 67448
rect 0 63928 800 64048
rect 99200 61208 100000 61328
rect 0 57808 800 57928
rect 99200 54408 100000 54528
rect 0 51008 800 51128
rect 99200 48288 100000 48408
rect 0 44888 800 45008
rect 99200 41488 100000 41608
rect 0 38088 800 38208
rect 99200 35368 100000 35488
rect 0 31968 800 32088
rect 99200 28568 100000 28688
rect 0 25168 800 25288
rect 99200 22448 100000 22568
rect 0 19048 800 19168
rect 99200 15648 100000 15768
rect 0 12248 800 12368
rect 99200 9528 100000 9648
rect 0 6128 800 6248
rect 99200 2728 100000 2848
<< obsm3 >>
rect 800 96768 99200 97409
rect 880 96488 99200 96768
rect 800 93368 99200 96488
rect 800 93088 99120 93368
rect 800 89968 99200 93088
rect 880 89688 99200 89968
rect 800 87248 99200 89688
rect 800 86968 99120 87248
rect 800 83848 99200 86968
rect 880 83568 99200 83848
rect 800 80448 99200 83568
rect 800 80168 99120 80448
rect 800 77048 99200 80168
rect 880 76768 99200 77048
rect 800 74328 99200 76768
rect 800 74048 99120 74328
rect 800 70928 99200 74048
rect 880 70648 99200 70928
rect 800 67528 99200 70648
rect 800 67248 99120 67528
rect 800 64128 99200 67248
rect 880 63848 99200 64128
rect 800 61408 99200 63848
rect 800 61128 99120 61408
rect 800 58008 99200 61128
rect 880 57728 99200 58008
rect 800 54608 99200 57728
rect 800 54328 99120 54608
rect 800 51208 99200 54328
rect 880 50928 99200 51208
rect 800 48488 99200 50928
rect 800 48208 99120 48488
rect 800 45088 99200 48208
rect 880 44808 99200 45088
rect 800 41688 99200 44808
rect 800 41408 99120 41688
rect 800 38288 99200 41408
rect 880 38008 99200 38288
rect 800 35568 99200 38008
rect 800 35288 99120 35568
rect 800 32168 99200 35288
rect 880 31888 99200 32168
rect 800 28768 99200 31888
rect 800 28488 99120 28768
rect 800 25368 99200 28488
rect 880 25088 99200 25368
rect 800 22648 99200 25088
rect 800 22368 99120 22648
rect 800 19248 99200 22368
rect 880 18968 99200 19248
rect 800 15848 99200 18968
rect 800 15568 99120 15848
rect 800 12448 99200 15568
rect 880 12168 99200 12448
rect 800 9728 99200 12168
rect 800 9448 99120 9728
rect 800 6328 99200 9448
rect 880 6048 99200 6328
rect 800 2928 99200 6048
rect 800 2648 99120 2928
rect 800 2143 99200 2648
<< metal4 >>
rect 4208 2128 4528 97424
rect 19568 2128 19888 97424
rect 34928 2128 35248 97424
rect 50288 2128 50608 97424
rect 65648 2128 65968 97424
rect 81008 2128 81328 97424
rect 96368 2128 96688 97424
<< obsm4 >>
rect 23795 2347 34848 97205
rect 35328 2347 50208 97205
rect 50688 2347 65568 97205
rect 66048 2347 80928 97205
rect 81408 2347 82373 97205
<< labels >>
rlabel metal3 s 0 12248 800 12368 6 io_msg[0]
port 1 nsew signal input
rlabel metal3 s 99200 35368 100000 35488 6 io_msg[10]
port 2 nsew signal input
rlabel metal3 s 99200 2728 100000 2848 6 io_msg[11]
port 3 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_msg[12]
port 4 nsew signal input
rlabel metal2 s 45098 99200 45154 100000 6 io_msg[13]
port 5 nsew signal input
rlabel metal2 s 20626 99200 20682 100000 6 io_msg[14]
port 6 nsew signal input
rlabel metal2 s 2594 99200 2650 100000 6 io_msg[15]
port 7 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 io_msg[16]
port 8 nsew signal input
rlabel metal3 s 99200 67328 100000 67448 6 io_msg[17]
port 9 nsew signal input
rlabel metal3 s 99200 15648 100000 15768 6 io_msg[18]
port 10 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 io_msg[19]
port 11 nsew signal input
rlabel metal2 s 39302 99200 39358 100000 6 io_msg[1]
port 12 nsew signal input
rlabel metal2 s 69570 99200 69626 100000 6 io_msg[20]
port 13 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 io_msg[21]
port 14 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 io_msg[22]
port 15 nsew signal input
rlabel metal3 s 99200 54408 100000 54528 6 io_msg[23]
port 16 nsew signal input
rlabel metal3 s 99200 28568 100000 28688 6 io_msg[24]
port 17 nsew signal input
rlabel metal2 s 57334 99200 57390 100000 6 io_msg[25]
port 18 nsew signal input
rlabel metal3 s 99200 87048 100000 87168 6 io_msg[26]
port 19 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 io_msg[27]
port 20 nsew signal input
rlabel metal3 s 99200 61208 100000 61328 6 io_msg[28]
port 21 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 io_msg[29]
port 22 nsew signal input
rlabel metal3 s 99200 93168 100000 93288 6 io_msg[2]
port 23 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 io_msg[30]
port 24 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 io_msg[31]
port 25 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 io_msg[3]
port 26 nsew signal input
rlabel metal2 s 8390 99200 8446 100000 6 io_msg[4]
port 27 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 io_msg[5]
port 28 nsew signal input
rlabel metal2 s 63774 99200 63830 100000 6 io_msg[6]
port 29 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 io_msg[7]
port 30 nsew signal input
rlabel metal3 s 99200 9528 100000 9648 6 io_msg[8]
port 31 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 io_msg[9]
port 32 nsew signal input
rlabel metal3 s 99200 22448 100000 22568 6 io_msg_out[0]
port 33 nsew signal output
rlabel metal2 s 81806 99200 81862 100000 6 io_msg_out[10]
port 34 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 io_msg_out[11]
port 35 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_msg_out[12]
port 36 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_msg_out[13]
port 37 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 io_msg_out[14]
port 38 nsew signal output
rlabel metal2 s 76010 99200 76066 100000 6 io_msg_out[15]
port 39 nsew signal output
rlabel metal2 s 94042 99200 94098 100000 6 io_msg_out[16]
port 40 nsew signal output
rlabel metal2 s 27066 99200 27122 100000 6 io_msg_out[17]
port 41 nsew signal output
rlabel metal2 s 51538 99200 51594 100000 6 io_msg_out[18]
port 42 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 io_msg_out[19]
port 43 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_msg_out[1]
port 44 nsew signal output
rlabel metal3 s 99200 80248 100000 80368 6 io_msg_out[20]
port 45 nsew signal output
rlabel metal2 s 99838 99200 99894 100000 6 io_msg_out[21]
port 46 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 io_msg_out[22]
port 47 nsew signal output
rlabel metal3 s 99200 74128 100000 74248 6 io_msg_out[23]
port 48 nsew signal output
rlabel metal2 s 97262 0 97318 800 6 io_msg_out[24]
port 49 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 io_msg_out[25]
port 50 nsew signal output
rlabel metal3 s 0 6128 800 6248 6 io_msg_out[26]
port 51 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 io_msg_out[27]
port 52 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 io_msg_out[28]
port 53 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 io_msg_out[29]
port 54 nsew signal output
rlabel metal3 s 99200 48288 100000 48408 6 io_msg_out[2]
port 55 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 io_msg_out[30]
port 56 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 io_msg_out[31]
port 57 nsew signal output
rlabel metal2 s 88246 99200 88302 100000 6 io_msg_out[3]
port 58 nsew signal output
rlabel metal2 s 14830 99200 14886 100000 6 io_msg_out[4]
port 59 nsew signal output
rlabel metal2 s 32862 99200 32918 100000 6 io_msg_out[5]
port 60 nsew signal output
rlabel metal2 s 66994 0 67050 800 6 io_msg_out[6]
port 61 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 io_msg_out[7]
port 62 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 io_msg_out[8]
port 63 nsew signal output
rlabel metal3 s 99200 41488 100000 41608 6 io_msg_out[9]
port 64 nsew signal output
rlabel metal4 s 4208 2128 4528 97424 6 vccd1
port 65 nsew power input
rlabel metal4 s 34928 2128 35248 97424 6 vccd1
port 65 nsew power input
rlabel metal4 s 65648 2128 65968 97424 6 vccd1
port 65 nsew power input
rlabel metal4 s 96368 2128 96688 97424 6 vccd1
port 65 nsew power input
rlabel metal4 s 19568 2128 19888 97424 6 vssd1
port 66 nsew ground input
rlabel metal4 s 50288 2128 50608 97424 6 vssd1
port 66 nsew ground input
rlabel metal4 s 81008 2128 81328 97424 6 vssd1
port 66 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12263502
string GDS_FILE /home/askartos/sandbox/caravel_tutorial/fossiAES/openlane/sbox/runs/sbox/results/finishing/sbox.magic.gds
string GDS_START 867496
<< end >>

