VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO aes
  CLASS BLOCK ;
  FOREIGN aes ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 800.000 ;
  PIN clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 796.000 93.750 800.000 ;
    END
  END clock
  PIN io_wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END io_wbs_ack_o
  PIN io_wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 646.040 800.000 646.640 ;
    END
  END io_wbs_adr_i[0]
  PIN io_wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END io_wbs_adr_i[10]
  PIN io_wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END io_wbs_adr_i[11]
  PIN io_wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 796.000 505.910 800.000 ;
    END
  END io_wbs_adr_i[12]
  PIN io_wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 796.000 592.850 800.000 ;
    END
  END io_wbs_adr_i[13]
  PIN io_wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END io_wbs_adr_i[14]
  PIN io_wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END io_wbs_adr_i[15]
  PIN io_wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 550.840 800.000 551.440 ;
    END
  END io_wbs_adr_i[16]
  PIN io_wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 428.440 800.000 429.040 ;
    END
  END io_wbs_adr_i[17]
  PIN io_wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 23.840 800.000 24.440 ;
    END
  END io_wbs_adr_i[18]
  PIN io_wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 622.240 4.000 622.840 ;
    END
  END io_wbs_adr_i[19]
  PIN io_wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END io_wbs_adr_i[1]
  PIN io_wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END io_wbs_adr_i[20]
  PIN io_wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 176.840 800.000 177.440 ;
    END
  END io_wbs_adr_i[21]
  PIN io_wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 796.000 418.970 800.000 ;
    END
  END io_wbs_adr_i[22]
  PIN io_wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END io_wbs_adr_i[23]
  PIN io_wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 796.000 241.870 800.000 ;
    END
  END io_wbs_adr_i[24]
  PIN io_wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 737.840 800.000 738.440 ;
    END
  END io_wbs_adr_i[25]
  PIN io_wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 796.000 476.930 800.000 ;
    END
  END io_wbs_adr_i[26]
  PIN io_wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 146.240 800.000 146.840 ;
    END
  END io_wbs_adr_i[27]
  PIN io_wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END io_wbs_adr_i[28]
  PIN io_wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END io_wbs_adr_i[29]
  PIN io_wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END io_wbs_adr_i[2]
  PIN io_wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 115.640 800.000 116.240 ;
    END
  END io_wbs_adr_i[30]
  PIN io_wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 796.000 563.870 800.000 ;
    END
  END io_wbs_adr_i[31]
  PIN io_wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END io_wbs_adr_i[3]
  PIN io_wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END io_wbs_adr_i[4]
  PIN io_wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END io_wbs_adr_i[5]
  PIN io_wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 796.000 740.970 800.000 ;
    END
  END io_wbs_adr_i[6]
  PIN io_wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END io_wbs_adr_i[7]
  PIN io_wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END io_wbs_adr_i[8]
  PIN io_wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 796.000 798.930 800.000 ;
    END
  END io_wbs_adr_i[9]
  PIN io_wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 796.000 654.030 800.000 ;
    END
  END io_wbs_cyc_i
  PIN io_wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 676.640 800.000 677.240 ;
    END
  END io_wbs_dat_i[0]
  PIN io_wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 768.440 800.000 769.040 ;
    END
  END io_wbs_dat_i[10]
  PIN io_wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 333.240 800.000 333.840 ;
    END
  END io_wbs_dat_i[11]
  PIN io_wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 272.040 800.000 272.640 ;
    END
  END io_wbs_dat_i[12]
  PIN io_wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 796.000 270.850 800.000 ;
    END
  END io_wbs_dat_i[13]
  PIN io_wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 796.000 299.830 800.000 ;
    END
  END io_wbs_dat_i[14]
  PIN io_wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 615.440 800.000 616.040 ;
    END
  END io_wbs_dat_i[15]
  PIN io_wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 796.000 386.770 800.000 ;
    END
  END io_wbs_dat_i[16]
  PIN io_wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END io_wbs_dat_i[17]
  PIN io_wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 796.000 328.810 800.000 ;
    END
  END io_wbs_dat_i[18]
  PIN io_wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 0.000 795.710 4.000 ;
    END
  END io_wbs_dat_i[19]
  PIN io_wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 796.000 447.950 800.000 ;
    END
  END io_wbs_dat_i[1]
  PIN io_wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END io_wbs_dat_i[20]
  PIN io_wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 796.000 209.670 800.000 ;
    END
  END io_wbs_dat_i[21]
  PIN io_wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 54.440 800.000 55.040 ;
    END
  END io_wbs_dat_i[22]
  PIN io_wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 707.240 800.000 707.840 ;
    END
  END io_wbs_dat_i[23]
  PIN io_wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 796.000 683.010 800.000 ;
    END
  END io_wbs_dat_i[24]
  PIN io_wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END io_wbs_dat_i[25]
  PIN io_wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END io_wbs_dat_i[26]
  PIN io_wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 210.840 800.000 211.440 ;
    END
  END io_wbs_dat_i[27]
  PIN io_wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_wbs_dat_i[28]
  PIN io_wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END io_wbs_dat_i[29]
  PIN io_wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END io_wbs_dat_i[2]
  PIN io_wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 796.000 151.710 800.000 ;
    END
  END io_wbs_dat_i[30]
  PIN io_wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END io_wbs_dat_i[31]
  PIN io_wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 744.640 4.000 745.240 ;
    END
  END io_wbs_dat_i[3]
  PIN io_wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_wbs_dat_i[4]
  PIN io_wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END io_wbs_dat_i[5]
  PIN io_wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END io_wbs_dat_i[6]
  PIN io_wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END io_wbs_dat_i[7]
  PIN io_wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 397.840 800.000 398.440 ;
    END
  END io_wbs_dat_i[8]
  PIN io_wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 241.440 800.000 242.040 ;
    END
  END io_wbs_dat_i[9]
  PIN io_wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END io_wbs_dat_o[0]
  PIN io_wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_wbs_dat_o[10]
  PIN io_wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END io_wbs_dat_o[11]
  PIN io_wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_wbs_dat_o[12]
  PIN io_wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 302.640 800.000 303.240 ;
    END
  END io_wbs_dat_o[13]
  PIN io_wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 520.240 800.000 520.840 ;
    END
  END io_wbs_dat_o[14]
  PIN io_wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END io_wbs_dat_o[15]
  PIN io_wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 581.440 800.000 582.040 ;
    END
  END io_wbs_dat_o[16]
  PIN io_wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END io_wbs_dat_o[17]
  PIN io_wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 796.000 3.590 800.000 ;
    END
  END io_wbs_dat_o[18]
  PIN io_wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END io_wbs_dat_o[19]
  PIN io_wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END io_wbs_dat_o[1]
  PIN io_wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END io_wbs_dat_o[20]
  PIN io_wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 796.000 122.730 800.000 ;
    END
  END io_wbs_dat_o[21]
  PIN io_wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 796.000 357.790 800.000 ;
    END
  END io_wbs_dat_o[22]
  PIN io_wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END io_wbs_dat_o[23]
  PIN io_wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.240 4.000 775.840 ;
    END
  END io_wbs_dat_o[24]
  PIN io_wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_wbs_dat_o[25]
  PIN io_wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END io_wbs_dat_o[26]
  PIN io_wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 796.000 711.990 800.000 ;
    END
  END io_wbs_dat_o[27]
  PIN io_wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 796.000 534.890 800.000 ;
    END
  END io_wbs_dat_o[28]
  PIN io_wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 0.000 351.350 4.000 ;
    END
  END io_wbs_dat_o[29]
  PIN io_wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 796.000 769.950 800.000 ;
    END
  END io_wbs_dat_o[2]
  PIN io_wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 85.040 800.000 85.640 ;
    END
  END io_wbs_dat_o[30]
  PIN io_wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 796.000 35.790 800.000 ;
    END
  END io_wbs_dat_o[31]
  PIN io_wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 459.040 800.000 459.640 ;
    END
  END io_wbs_dat_o[3]
  PIN io_wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END io_wbs_dat_o[4]
  PIN io_wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END io_wbs_dat_o[5]
  PIN io_wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END io_wbs_dat_o[6]
  PIN io_wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 489.640 800.000 490.240 ;
    END
  END io_wbs_dat_o[7]
  PIN io_wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END io_wbs_dat_o[8]
  PIN io_wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_wbs_dat_o[9]
  PIN io_wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 796.000 625.050 800.000 ;
    END
  END io_wbs_sel_i[0]
  PIN io_wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 796.000 64.770 800.000 ;
    END
  END io_wbs_sel_i[1]
  PIN io_wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 796.000 180.690 800.000 ;
    END
  END io_wbs_sel_i[2]
  PIN io_wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END io_wbs_sel_i[3]
  PIN io_wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END io_wbs_stb_i
  PIN io_wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 714.040 4.000 714.640 ;
    END
  END io_wbs_we_i
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.000 363.840 800.000 364.440 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 794.420 788.885 ;
      LAYER met1 ;
        RECT 0.070 10.640 795.730 789.440 ;
      LAYER met2 ;
        RECT 0.100 795.720 3.030 796.690 ;
        RECT 3.870 795.720 35.230 796.690 ;
        RECT 36.070 795.720 64.210 796.690 ;
        RECT 65.050 795.720 93.190 796.690 ;
        RECT 94.030 795.720 122.170 796.690 ;
        RECT 123.010 795.720 151.150 796.690 ;
        RECT 151.990 795.720 180.130 796.690 ;
        RECT 180.970 795.720 209.110 796.690 ;
        RECT 209.950 795.720 241.310 796.690 ;
        RECT 242.150 795.720 270.290 796.690 ;
        RECT 271.130 795.720 299.270 796.690 ;
        RECT 300.110 795.720 328.250 796.690 ;
        RECT 329.090 795.720 357.230 796.690 ;
        RECT 358.070 795.720 386.210 796.690 ;
        RECT 387.050 795.720 418.410 796.690 ;
        RECT 419.250 795.720 447.390 796.690 ;
        RECT 448.230 795.720 476.370 796.690 ;
        RECT 477.210 795.720 505.350 796.690 ;
        RECT 506.190 795.720 534.330 796.690 ;
        RECT 535.170 795.720 563.310 796.690 ;
        RECT 564.150 795.720 592.290 796.690 ;
        RECT 593.130 795.720 624.490 796.690 ;
        RECT 625.330 795.720 653.470 796.690 ;
        RECT 654.310 795.720 682.450 796.690 ;
        RECT 683.290 795.720 711.430 796.690 ;
        RECT 712.270 795.720 740.410 796.690 ;
        RECT 741.250 795.720 769.390 796.690 ;
        RECT 770.230 795.720 795.700 796.690 ;
        RECT 0.100 4.280 795.700 795.720 ;
        RECT 0.650 4.000 28.790 4.280 ;
        RECT 29.630 4.000 57.770 4.280 ;
        RECT 58.610 4.000 86.750 4.280 ;
        RECT 87.590 4.000 115.730 4.280 ;
        RECT 116.570 4.000 144.710 4.280 ;
        RECT 145.550 4.000 173.690 4.280 ;
        RECT 174.530 4.000 205.890 4.280 ;
        RECT 206.730 4.000 234.870 4.280 ;
        RECT 235.710 4.000 263.850 4.280 ;
        RECT 264.690 4.000 292.830 4.280 ;
        RECT 293.670 4.000 321.810 4.280 ;
        RECT 322.650 4.000 350.790 4.280 ;
        RECT 351.630 4.000 379.770 4.280 ;
        RECT 380.610 4.000 411.970 4.280 ;
        RECT 412.810 4.000 440.950 4.280 ;
        RECT 441.790 4.000 469.930 4.280 ;
        RECT 470.770 4.000 498.910 4.280 ;
        RECT 499.750 4.000 527.890 4.280 ;
        RECT 528.730 4.000 556.870 4.280 ;
        RECT 557.710 4.000 589.070 4.280 ;
        RECT 589.910 4.000 618.050 4.280 ;
        RECT 618.890 4.000 647.030 4.280 ;
        RECT 647.870 4.000 676.010 4.280 ;
        RECT 676.850 4.000 704.990 4.280 ;
        RECT 705.830 4.000 733.970 4.280 ;
        RECT 734.810 4.000 762.950 4.280 ;
        RECT 763.790 4.000 795.150 4.280 ;
      LAYER met3 ;
        RECT 4.000 776.240 796.000 788.965 ;
        RECT 4.400 774.840 796.000 776.240 ;
        RECT 4.000 769.440 796.000 774.840 ;
        RECT 4.000 768.040 795.600 769.440 ;
        RECT 4.000 745.640 796.000 768.040 ;
        RECT 4.400 744.240 796.000 745.640 ;
        RECT 4.000 738.840 796.000 744.240 ;
        RECT 4.000 737.440 795.600 738.840 ;
        RECT 4.000 715.040 796.000 737.440 ;
        RECT 4.400 713.640 796.000 715.040 ;
        RECT 4.000 708.240 796.000 713.640 ;
        RECT 4.000 706.840 795.600 708.240 ;
        RECT 4.000 684.440 796.000 706.840 ;
        RECT 4.400 683.040 796.000 684.440 ;
        RECT 4.000 677.640 796.000 683.040 ;
        RECT 4.000 676.240 795.600 677.640 ;
        RECT 4.000 653.840 796.000 676.240 ;
        RECT 4.400 652.440 796.000 653.840 ;
        RECT 4.000 647.040 796.000 652.440 ;
        RECT 4.000 645.640 795.600 647.040 ;
        RECT 4.000 623.240 796.000 645.640 ;
        RECT 4.400 621.840 796.000 623.240 ;
        RECT 4.000 616.440 796.000 621.840 ;
        RECT 4.000 615.040 795.600 616.440 ;
        RECT 4.000 589.240 796.000 615.040 ;
        RECT 4.400 587.840 796.000 589.240 ;
        RECT 4.000 582.440 796.000 587.840 ;
        RECT 4.000 581.040 795.600 582.440 ;
        RECT 4.000 558.640 796.000 581.040 ;
        RECT 4.400 557.240 796.000 558.640 ;
        RECT 4.000 551.840 796.000 557.240 ;
        RECT 4.000 550.440 795.600 551.840 ;
        RECT 4.000 528.040 796.000 550.440 ;
        RECT 4.400 526.640 796.000 528.040 ;
        RECT 4.000 521.240 796.000 526.640 ;
        RECT 4.000 519.840 795.600 521.240 ;
        RECT 4.000 497.440 796.000 519.840 ;
        RECT 4.400 496.040 796.000 497.440 ;
        RECT 4.000 490.640 796.000 496.040 ;
        RECT 4.000 489.240 795.600 490.640 ;
        RECT 4.000 466.840 796.000 489.240 ;
        RECT 4.400 465.440 796.000 466.840 ;
        RECT 4.000 460.040 796.000 465.440 ;
        RECT 4.000 458.640 795.600 460.040 ;
        RECT 4.000 436.240 796.000 458.640 ;
        RECT 4.400 434.840 796.000 436.240 ;
        RECT 4.000 429.440 796.000 434.840 ;
        RECT 4.000 428.040 795.600 429.440 ;
        RECT 4.000 402.240 796.000 428.040 ;
        RECT 4.400 400.840 796.000 402.240 ;
        RECT 4.000 398.840 796.000 400.840 ;
        RECT 4.000 397.440 795.600 398.840 ;
        RECT 4.000 371.640 796.000 397.440 ;
        RECT 4.400 370.240 796.000 371.640 ;
        RECT 4.000 364.840 796.000 370.240 ;
        RECT 4.000 363.440 795.600 364.840 ;
        RECT 4.000 341.040 796.000 363.440 ;
        RECT 4.400 339.640 796.000 341.040 ;
        RECT 4.000 334.240 796.000 339.640 ;
        RECT 4.000 332.840 795.600 334.240 ;
        RECT 4.000 310.440 796.000 332.840 ;
        RECT 4.400 309.040 796.000 310.440 ;
        RECT 4.000 303.640 796.000 309.040 ;
        RECT 4.000 302.240 795.600 303.640 ;
        RECT 4.000 279.840 796.000 302.240 ;
        RECT 4.400 278.440 796.000 279.840 ;
        RECT 4.000 273.040 796.000 278.440 ;
        RECT 4.000 271.640 795.600 273.040 ;
        RECT 4.000 249.240 796.000 271.640 ;
        RECT 4.400 247.840 796.000 249.240 ;
        RECT 4.000 242.440 796.000 247.840 ;
        RECT 4.000 241.040 795.600 242.440 ;
        RECT 4.000 218.640 796.000 241.040 ;
        RECT 4.400 217.240 796.000 218.640 ;
        RECT 4.000 211.840 796.000 217.240 ;
        RECT 4.000 210.440 795.600 211.840 ;
        RECT 4.000 184.640 796.000 210.440 ;
        RECT 4.400 183.240 796.000 184.640 ;
        RECT 4.000 177.840 796.000 183.240 ;
        RECT 4.000 176.440 795.600 177.840 ;
        RECT 4.000 154.040 796.000 176.440 ;
        RECT 4.400 152.640 796.000 154.040 ;
        RECT 4.000 147.240 796.000 152.640 ;
        RECT 4.000 145.840 795.600 147.240 ;
        RECT 4.000 123.440 796.000 145.840 ;
        RECT 4.400 122.040 796.000 123.440 ;
        RECT 4.000 116.640 796.000 122.040 ;
        RECT 4.000 115.240 795.600 116.640 ;
        RECT 4.000 92.840 796.000 115.240 ;
        RECT 4.400 91.440 796.000 92.840 ;
        RECT 4.000 86.040 796.000 91.440 ;
        RECT 4.000 84.640 795.600 86.040 ;
        RECT 4.000 62.240 796.000 84.640 ;
        RECT 4.400 60.840 796.000 62.240 ;
        RECT 4.000 55.440 796.000 60.840 ;
        RECT 4.000 54.040 795.600 55.440 ;
        RECT 4.000 31.640 796.000 54.040 ;
        RECT 4.400 30.240 796.000 31.640 ;
        RECT 4.000 24.840 796.000 30.240 ;
        RECT 4.000 23.440 795.600 24.840 ;
        RECT 4.000 10.715 796.000 23.440 ;
      LAYER met4 ;
        RECT 101.495 44.375 174.240 787.945 ;
        RECT 176.640 44.375 251.040 787.945 ;
        RECT 253.440 44.375 327.840 787.945 ;
        RECT 330.240 44.375 404.640 787.945 ;
        RECT 407.040 44.375 481.440 787.945 ;
        RECT 483.840 44.375 558.240 787.945 ;
        RECT 560.640 44.375 635.040 787.945 ;
        RECT 637.440 44.375 669.465 787.945 ;
  END
END aes
END LIBRARY

