module sbox(
  input  [31:0] io_msg,
  output [31:0] io_msg_out
);
  wire [7:0] _GEN_1 = 8'h1 == io_msg[7:0] ? 8'h7c : 8'h63; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_2 = 8'h2 == io_msg[7:0] ? 8'h77 : _GEN_1; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_3 = 8'h3 == io_msg[7:0] ? 8'h7b : _GEN_2; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_4 = 8'h4 == io_msg[7:0] ? 8'hf2 : _GEN_3; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_5 = 8'h5 == io_msg[7:0] ? 8'h6b : _GEN_4; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_6 = 8'h6 == io_msg[7:0] ? 8'h6f : _GEN_5; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_7 = 8'h7 == io_msg[7:0] ? 8'hc5 : _GEN_6; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_8 = 8'h8 == io_msg[7:0] ? 8'h30 : _GEN_7; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_9 = 8'h9 == io_msg[7:0] ? 8'h1 : _GEN_8; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_10 = 8'ha == io_msg[7:0] ? 8'h67 : _GEN_9; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_11 = 8'hb == io_msg[7:0] ? 8'h2b : _GEN_10; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_12 = 8'hc == io_msg[7:0] ? 8'hfe : _GEN_11; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_13 = 8'hd == io_msg[7:0] ? 8'hd7 : _GEN_12; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_14 = 8'he == io_msg[7:0] ? 8'hab : _GEN_13; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_15 = 8'hf == io_msg[7:0] ? 8'h76 : _GEN_14; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_16 = 8'h10 == io_msg[7:0] ? 8'hca : _GEN_15; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_17 = 8'h11 == io_msg[7:0] ? 8'h82 : _GEN_16; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_18 = 8'h12 == io_msg[7:0] ? 8'hc9 : _GEN_17; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_19 = 8'h13 == io_msg[7:0] ? 8'h7d : _GEN_18; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_20 = 8'h14 == io_msg[7:0] ? 8'hfa : _GEN_19; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_21 = 8'h15 == io_msg[7:0] ? 8'h59 : _GEN_20; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_22 = 8'h16 == io_msg[7:0] ? 8'h47 : _GEN_21; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_23 = 8'h17 == io_msg[7:0] ? 8'hf0 : _GEN_22; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_24 = 8'h18 == io_msg[7:0] ? 8'had : _GEN_23; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_25 = 8'h19 == io_msg[7:0] ? 8'hd4 : _GEN_24; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_26 = 8'h1a == io_msg[7:0] ? 8'ha2 : _GEN_25; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_27 = 8'h1b == io_msg[7:0] ? 8'haf : _GEN_26; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_28 = 8'h1c == io_msg[7:0] ? 8'h9c : _GEN_27; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_29 = 8'h1d == io_msg[7:0] ? 8'ha4 : _GEN_28; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_30 = 8'h1e == io_msg[7:0] ? 8'h72 : _GEN_29; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_31 = 8'h1f == io_msg[7:0] ? 8'hc0 : _GEN_30; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_32 = 8'h20 == io_msg[7:0] ? 8'hb7 : _GEN_31; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_33 = 8'h21 == io_msg[7:0] ? 8'hfd : _GEN_32; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_34 = 8'h22 == io_msg[7:0] ? 8'h93 : _GEN_33; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_35 = 8'h23 == io_msg[7:0] ? 8'h26 : _GEN_34; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_36 = 8'h24 == io_msg[7:0] ? 8'h36 : _GEN_35; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_37 = 8'h25 == io_msg[7:0] ? 8'h3f : _GEN_36; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_38 = 8'h26 == io_msg[7:0] ? 8'hf7 : _GEN_37; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_39 = 8'h27 == io_msg[7:0] ? 8'hcc : _GEN_38; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_40 = 8'h28 == io_msg[7:0] ? 8'h34 : _GEN_39; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_41 = 8'h29 == io_msg[7:0] ? 8'ha5 : _GEN_40; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_42 = 8'h2a == io_msg[7:0] ? 8'he5 : _GEN_41; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_43 = 8'h2b == io_msg[7:0] ? 8'hf1 : _GEN_42; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_44 = 8'h2c == io_msg[7:0] ? 8'h71 : _GEN_43; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_45 = 8'h2d == io_msg[7:0] ? 8'hd8 : _GEN_44; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_46 = 8'h2e == io_msg[7:0] ? 8'h31 : _GEN_45; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_47 = 8'h2f == io_msg[7:0] ? 8'h15 : _GEN_46; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_48 = 8'h30 == io_msg[7:0] ? 8'h4 : _GEN_47; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_49 = 8'h31 == io_msg[7:0] ? 8'hc7 : _GEN_48; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_50 = 8'h32 == io_msg[7:0] ? 8'h23 : _GEN_49; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_51 = 8'h33 == io_msg[7:0] ? 8'hc3 : _GEN_50; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_52 = 8'h34 == io_msg[7:0] ? 8'h18 : _GEN_51; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_53 = 8'h35 == io_msg[7:0] ? 8'h96 : _GEN_52; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_54 = 8'h36 == io_msg[7:0] ? 8'h5 : _GEN_53; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_55 = 8'h37 == io_msg[7:0] ? 8'h9a : _GEN_54; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_56 = 8'h38 == io_msg[7:0] ? 8'h7 : _GEN_55; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_57 = 8'h39 == io_msg[7:0] ? 8'h12 : _GEN_56; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_58 = 8'h3a == io_msg[7:0] ? 8'h80 : _GEN_57; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_59 = 8'h3b == io_msg[7:0] ? 8'he2 : _GEN_58; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_60 = 8'h3c == io_msg[7:0] ? 8'heb : _GEN_59; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_61 = 8'h3d == io_msg[7:0] ? 8'h27 : _GEN_60; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_62 = 8'h3e == io_msg[7:0] ? 8'hb2 : _GEN_61; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_63 = 8'h3f == io_msg[7:0] ? 8'h75 : _GEN_62; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_64 = 8'h40 == io_msg[7:0] ? 8'h9 : _GEN_63; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_65 = 8'h41 == io_msg[7:0] ? 8'h83 : _GEN_64; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_66 = 8'h42 == io_msg[7:0] ? 8'h2c : _GEN_65; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_67 = 8'h43 == io_msg[7:0] ? 8'h1a : _GEN_66; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_68 = 8'h44 == io_msg[7:0] ? 8'h1b : _GEN_67; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_69 = 8'h45 == io_msg[7:0] ? 8'h6e : _GEN_68; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_70 = 8'h46 == io_msg[7:0] ? 8'h5a : _GEN_69; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_71 = 8'h47 == io_msg[7:0] ? 8'ha0 : _GEN_70; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_72 = 8'h48 == io_msg[7:0] ? 8'h52 : _GEN_71; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_73 = 8'h49 == io_msg[7:0] ? 8'h3b : _GEN_72; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_74 = 8'h4a == io_msg[7:0] ? 8'hd6 : _GEN_73; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_75 = 8'h4b == io_msg[7:0] ? 8'hb3 : _GEN_74; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_76 = 8'h4c == io_msg[7:0] ? 8'h29 : _GEN_75; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_77 = 8'h4d == io_msg[7:0] ? 8'he3 : _GEN_76; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_78 = 8'h4e == io_msg[7:0] ? 8'h2f : _GEN_77; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_79 = 8'h4f == io_msg[7:0] ? 8'h84 : _GEN_78; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_80 = 8'h50 == io_msg[7:0] ? 8'h53 : _GEN_79; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_81 = 8'h51 == io_msg[7:0] ? 8'hd1 : _GEN_80; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_82 = 8'h52 == io_msg[7:0] ? 8'h0 : _GEN_81; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_83 = 8'h53 == io_msg[7:0] ? 8'hed : _GEN_82; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_84 = 8'h54 == io_msg[7:0] ? 8'h20 : _GEN_83; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_85 = 8'h55 == io_msg[7:0] ? 8'hfc : _GEN_84; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_86 = 8'h56 == io_msg[7:0] ? 8'hb1 : _GEN_85; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_87 = 8'h57 == io_msg[7:0] ? 8'h5b : _GEN_86; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_88 = 8'h58 == io_msg[7:0] ? 8'h6a : _GEN_87; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_89 = 8'h59 == io_msg[7:0] ? 8'hcb : _GEN_88; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_90 = 8'h5a == io_msg[7:0] ? 8'hbe : _GEN_89; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_91 = 8'h5b == io_msg[7:0] ? 8'h39 : _GEN_90; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_92 = 8'h5c == io_msg[7:0] ? 8'h4a : _GEN_91; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_93 = 8'h5d == io_msg[7:0] ? 8'h4c : _GEN_92; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_94 = 8'h5e == io_msg[7:0] ? 8'h58 : _GEN_93; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_95 = 8'h5f == io_msg[7:0] ? 8'hcf : _GEN_94; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_96 = 8'h60 == io_msg[7:0] ? 8'hd0 : _GEN_95; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_97 = 8'h61 == io_msg[7:0] ? 8'hef : _GEN_96; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_98 = 8'h62 == io_msg[7:0] ? 8'haa : _GEN_97; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_99 = 8'h63 == io_msg[7:0] ? 8'hfb : _GEN_98; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_100 = 8'h64 == io_msg[7:0] ? 8'h43 : _GEN_99; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_101 = 8'h65 == io_msg[7:0] ? 8'h4d : _GEN_100; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_102 = 8'h66 == io_msg[7:0] ? 8'h33 : _GEN_101; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_103 = 8'h67 == io_msg[7:0] ? 8'h85 : _GEN_102; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_104 = 8'h68 == io_msg[7:0] ? 8'h45 : _GEN_103; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_105 = 8'h69 == io_msg[7:0] ? 8'hf9 : _GEN_104; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_106 = 8'h6a == io_msg[7:0] ? 8'h2 : _GEN_105; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_107 = 8'h6b == io_msg[7:0] ? 8'h7f : _GEN_106; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_108 = 8'h6c == io_msg[7:0] ? 8'h50 : _GEN_107; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_109 = 8'h6d == io_msg[7:0] ? 8'h3c : _GEN_108; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_110 = 8'h6e == io_msg[7:0] ? 8'h9f : _GEN_109; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_111 = 8'h6f == io_msg[7:0] ? 8'ha8 : _GEN_110; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_112 = 8'h70 == io_msg[7:0] ? 8'h51 : _GEN_111; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_113 = 8'h71 == io_msg[7:0] ? 8'ha3 : _GEN_112; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_114 = 8'h72 == io_msg[7:0] ? 8'h40 : _GEN_113; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_115 = 8'h73 == io_msg[7:0] ? 8'h8f : _GEN_114; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_116 = 8'h74 == io_msg[7:0] ? 8'h92 : _GEN_115; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_117 = 8'h75 == io_msg[7:0] ? 8'h9d : _GEN_116; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_118 = 8'h76 == io_msg[7:0] ? 8'h38 : _GEN_117; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_119 = 8'h77 == io_msg[7:0] ? 8'hf5 : _GEN_118; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_120 = 8'h78 == io_msg[7:0] ? 8'hbc : _GEN_119; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_121 = 8'h79 == io_msg[7:0] ? 8'hb6 : _GEN_120; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_122 = 8'h7a == io_msg[7:0] ? 8'hda : _GEN_121; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_123 = 8'h7b == io_msg[7:0] ? 8'h21 : _GEN_122; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_124 = 8'h7c == io_msg[7:0] ? 8'h10 : _GEN_123; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_125 = 8'h7d == io_msg[7:0] ? 8'hff : _GEN_124; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_126 = 8'h7e == io_msg[7:0] ? 8'hf3 : _GEN_125; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_127 = 8'h7f == io_msg[7:0] ? 8'hd2 : _GEN_126; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_128 = 8'h80 == io_msg[7:0] ? 8'hcd : _GEN_127; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_129 = 8'h81 == io_msg[7:0] ? 8'hc : _GEN_128; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_130 = 8'h82 == io_msg[7:0] ? 8'h13 : _GEN_129; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_131 = 8'h83 == io_msg[7:0] ? 8'hec : _GEN_130; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_132 = 8'h84 == io_msg[7:0] ? 8'h5f : _GEN_131; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_133 = 8'h85 == io_msg[7:0] ? 8'h97 : _GEN_132; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_134 = 8'h86 == io_msg[7:0] ? 8'h44 : _GEN_133; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_135 = 8'h87 == io_msg[7:0] ? 8'h17 : _GEN_134; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_136 = 8'h88 == io_msg[7:0] ? 8'hc4 : _GEN_135; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_137 = 8'h89 == io_msg[7:0] ? 8'ha7 : _GEN_136; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_138 = 8'h8a == io_msg[7:0] ? 8'h7e : _GEN_137; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_139 = 8'h8b == io_msg[7:0] ? 8'h3d : _GEN_138; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_140 = 8'h8c == io_msg[7:0] ? 8'h64 : _GEN_139; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_141 = 8'h8d == io_msg[7:0] ? 8'h5d : _GEN_140; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_142 = 8'h8e == io_msg[7:0] ? 8'h19 : _GEN_141; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_143 = 8'h8f == io_msg[7:0] ? 8'h73 : _GEN_142; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_144 = 8'h90 == io_msg[7:0] ? 8'h60 : _GEN_143; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_145 = 8'h91 == io_msg[7:0] ? 8'h81 : _GEN_144; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_146 = 8'h92 == io_msg[7:0] ? 8'h4f : _GEN_145; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_147 = 8'h93 == io_msg[7:0] ? 8'hdc : _GEN_146; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_148 = 8'h94 == io_msg[7:0] ? 8'h22 : _GEN_147; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_149 = 8'h95 == io_msg[7:0] ? 8'h2a : _GEN_148; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_150 = 8'h96 == io_msg[7:0] ? 8'h90 : _GEN_149; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_151 = 8'h97 == io_msg[7:0] ? 8'h88 : _GEN_150; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_152 = 8'h98 == io_msg[7:0] ? 8'h46 : _GEN_151; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_153 = 8'h99 == io_msg[7:0] ? 8'hee : _GEN_152; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_154 = 8'h9a == io_msg[7:0] ? 8'hb8 : _GEN_153; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_155 = 8'h9b == io_msg[7:0] ? 8'h14 : _GEN_154; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_156 = 8'h9c == io_msg[7:0] ? 8'hde : _GEN_155; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_157 = 8'h9d == io_msg[7:0] ? 8'h5e : _GEN_156; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_158 = 8'h9e == io_msg[7:0] ? 8'hb : _GEN_157; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_159 = 8'h9f == io_msg[7:0] ? 8'hdb : _GEN_158; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_160 = 8'ha0 == io_msg[7:0] ? 8'he0 : _GEN_159; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_161 = 8'ha1 == io_msg[7:0] ? 8'h32 : _GEN_160; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_162 = 8'ha2 == io_msg[7:0] ? 8'h3a : _GEN_161; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_163 = 8'ha3 == io_msg[7:0] ? 8'ha : _GEN_162; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_164 = 8'ha4 == io_msg[7:0] ? 8'h49 : _GEN_163; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_165 = 8'ha5 == io_msg[7:0] ? 8'h6 : _GEN_164; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_166 = 8'ha6 == io_msg[7:0] ? 8'h24 : _GEN_165; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_167 = 8'ha7 == io_msg[7:0] ? 8'h5c : _GEN_166; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_168 = 8'ha8 == io_msg[7:0] ? 8'hc2 : _GEN_167; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_169 = 8'ha9 == io_msg[7:0] ? 8'hd3 : _GEN_168; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_170 = 8'haa == io_msg[7:0] ? 8'hac : _GEN_169; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_171 = 8'hab == io_msg[7:0] ? 8'h62 : _GEN_170; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_172 = 8'hac == io_msg[7:0] ? 8'h91 : _GEN_171; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_173 = 8'had == io_msg[7:0] ? 8'h95 : _GEN_172; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_174 = 8'hae == io_msg[7:0] ? 8'he4 : _GEN_173; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_175 = 8'haf == io_msg[7:0] ? 8'h79 : _GEN_174; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_176 = 8'hb0 == io_msg[7:0] ? 8'he7 : _GEN_175; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_177 = 8'hb1 == io_msg[7:0] ? 8'hc8 : _GEN_176; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_178 = 8'hb2 == io_msg[7:0] ? 8'h37 : _GEN_177; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_179 = 8'hb3 == io_msg[7:0] ? 8'h6d : _GEN_178; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_180 = 8'hb4 == io_msg[7:0] ? 8'h8d : _GEN_179; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_181 = 8'hb5 == io_msg[7:0] ? 8'hd5 : _GEN_180; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_182 = 8'hb6 == io_msg[7:0] ? 8'h4e : _GEN_181; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_183 = 8'hb7 == io_msg[7:0] ? 8'ha9 : _GEN_182; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_184 = 8'hb8 == io_msg[7:0] ? 8'h6c : _GEN_183; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_185 = 8'hb9 == io_msg[7:0] ? 8'h56 : _GEN_184; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_186 = 8'hba == io_msg[7:0] ? 8'hf4 : _GEN_185; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_187 = 8'hbb == io_msg[7:0] ? 8'hea : _GEN_186; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_188 = 8'hbc == io_msg[7:0] ? 8'h65 : _GEN_187; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_189 = 8'hbd == io_msg[7:0] ? 8'h7a : _GEN_188; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_190 = 8'hbe == io_msg[7:0] ? 8'hae : _GEN_189; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_191 = 8'hbf == io_msg[7:0] ? 8'h8 : _GEN_190; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_192 = 8'hc0 == io_msg[7:0] ? 8'hba : _GEN_191; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_193 = 8'hc1 == io_msg[7:0] ? 8'h78 : _GEN_192; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_194 = 8'hc2 == io_msg[7:0] ? 8'h25 : _GEN_193; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_195 = 8'hc3 == io_msg[7:0] ? 8'h2e : _GEN_194; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_196 = 8'hc4 == io_msg[7:0] ? 8'h1c : _GEN_195; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_197 = 8'hc5 == io_msg[7:0] ? 8'ha6 : _GEN_196; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_198 = 8'hc6 == io_msg[7:0] ? 8'hb4 : _GEN_197; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_199 = 8'hc7 == io_msg[7:0] ? 8'hc6 : _GEN_198; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_200 = 8'hc8 == io_msg[7:0] ? 8'he8 : _GEN_199; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_201 = 8'hc9 == io_msg[7:0] ? 8'hdd : _GEN_200; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_202 = 8'hca == io_msg[7:0] ? 8'h74 : _GEN_201; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_203 = 8'hcb == io_msg[7:0] ? 8'h1f : _GEN_202; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_204 = 8'hcc == io_msg[7:0] ? 8'h4b : _GEN_203; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_205 = 8'hcd == io_msg[7:0] ? 8'hbd : _GEN_204; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_206 = 8'hce == io_msg[7:0] ? 8'h8b : _GEN_205; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_207 = 8'hcf == io_msg[7:0] ? 8'h8a : _GEN_206; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_208 = 8'hd0 == io_msg[7:0] ? 8'h70 : _GEN_207; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_209 = 8'hd1 == io_msg[7:0] ? 8'h3e : _GEN_208; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_210 = 8'hd2 == io_msg[7:0] ? 8'hb5 : _GEN_209; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_211 = 8'hd3 == io_msg[7:0] ? 8'h66 : _GEN_210; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_212 = 8'hd4 == io_msg[7:0] ? 8'h48 : _GEN_211; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_213 = 8'hd5 == io_msg[7:0] ? 8'h3 : _GEN_212; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_214 = 8'hd6 == io_msg[7:0] ? 8'hf6 : _GEN_213; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_215 = 8'hd7 == io_msg[7:0] ? 8'he : _GEN_214; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_216 = 8'hd8 == io_msg[7:0] ? 8'h61 : _GEN_215; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_217 = 8'hd9 == io_msg[7:0] ? 8'h35 : _GEN_216; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_218 = 8'hda == io_msg[7:0] ? 8'h57 : _GEN_217; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_219 = 8'hdb == io_msg[7:0] ? 8'hb9 : _GEN_218; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_220 = 8'hdc == io_msg[7:0] ? 8'h86 : _GEN_219; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_221 = 8'hdd == io_msg[7:0] ? 8'hc1 : _GEN_220; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_222 = 8'hde == io_msg[7:0] ? 8'h1d : _GEN_221; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_223 = 8'hdf == io_msg[7:0] ? 8'h9e : _GEN_222; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_224 = 8'he0 == io_msg[7:0] ? 8'he1 : _GEN_223; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_225 = 8'he1 == io_msg[7:0] ? 8'hf8 : _GEN_224; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_226 = 8'he2 == io_msg[7:0] ? 8'h98 : _GEN_225; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_227 = 8'he3 == io_msg[7:0] ? 8'h11 : _GEN_226; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_228 = 8'he4 == io_msg[7:0] ? 8'h69 : _GEN_227; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_229 = 8'he5 == io_msg[7:0] ? 8'hd9 : _GEN_228; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_230 = 8'he6 == io_msg[7:0] ? 8'h8e : _GEN_229; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_231 = 8'he7 == io_msg[7:0] ? 8'h94 : _GEN_230; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_232 = 8'he8 == io_msg[7:0] ? 8'h9b : _GEN_231; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_233 = 8'he9 == io_msg[7:0] ? 8'h1e : _GEN_232; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_234 = 8'hea == io_msg[7:0] ? 8'h87 : _GEN_233; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_235 = 8'heb == io_msg[7:0] ? 8'he9 : _GEN_234; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_236 = 8'hec == io_msg[7:0] ? 8'hce : _GEN_235; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_237 = 8'hed == io_msg[7:0] ? 8'h55 : _GEN_236; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_238 = 8'hee == io_msg[7:0] ? 8'h28 : _GEN_237; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_239 = 8'hef == io_msg[7:0] ? 8'hdf : _GEN_238; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_240 = 8'hf0 == io_msg[7:0] ? 8'h8c : _GEN_239; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_241 = 8'hf1 == io_msg[7:0] ? 8'ha1 : _GEN_240; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_242 = 8'hf2 == io_msg[7:0] ? 8'h89 : _GEN_241; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_243 = 8'hf3 == io_msg[7:0] ? 8'hd : _GEN_242; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_244 = 8'hf4 == io_msg[7:0] ? 8'hbf : _GEN_243; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_245 = 8'hf5 == io_msg[7:0] ? 8'he6 : _GEN_244; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_246 = 8'hf6 == io_msg[7:0] ? 8'h42 : _GEN_245; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_247 = 8'hf7 == io_msg[7:0] ? 8'h68 : _GEN_246; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_248 = 8'hf8 == io_msg[7:0] ? 8'h41 : _GEN_247; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_249 = 8'hf9 == io_msg[7:0] ? 8'h99 : _GEN_248; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_250 = 8'hfa == io_msg[7:0] ? 8'h2d : _GEN_249; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_251 = 8'hfb == io_msg[7:0] ? 8'hf : _GEN_250; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_252 = 8'hfc == io_msg[7:0] ? 8'hb0 : _GEN_251; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_253 = 8'hfd == io_msg[7:0] ? 8'h54 : _GEN_252; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_254 = 8'hfe == io_msg[7:0] ? 8'hbb : _GEN_253; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] sbox_out_0 = 8'hff == io_msg[7:0] ? 8'h16 : _GEN_254; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_257 = 8'h1 == io_msg[15:8] ? 8'h7c : 8'h63; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_258 = 8'h2 == io_msg[15:8] ? 8'h77 : _GEN_257; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_259 = 8'h3 == io_msg[15:8] ? 8'h7b : _GEN_258; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_260 = 8'h4 == io_msg[15:8] ? 8'hf2 : _GEN_259; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_261 = 8'h5 == io_msg[15:8] ? 8'h6b : _GEN_260; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_262 = 8'h6 == io_msg[15:8] ? 8'h6f : _GEN_261; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_263 = 8'h7 == io_msg[15:8] ? 8'hc5 : _GEN_262; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_264 = 8'h8 == io_msg[15:8] ? 8'h30 : _GEN_263; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_265 = 8'h9 == io_msg[15:8] ? 8'h1 : _GEN_264; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_266 = 8'ha == io_msg[15:8] ? 8'h67 : _GEN_265; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_267 = 8'hb == io_msg[15:8] ? 8'h2b : _GEN_266; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_268 = 8'hc == io_msg[15:8] ? 8'hfe : _GEN_267; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_269 = 8'hd == io_msg[15:8] ? 8'hd7 : _GEN_268; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_270 = 8'he == io_msg[15:8] ? 8'hab : _GEN_269; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_271 = 8'hf == io_msg[15:8] ? 8'h76 : _GEN_270; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_272 = 8'h10 == io_msg[15:8] ? 8'hca : _GEN_271; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_273 = 8'h11 == io_msg[15:8] ? 8'h82 : _GEN_272; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_274 = 8'h12 == io_msg[15:8] ? 8'hc9 : _GEN_273; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_275 = 8'h13 == io_msg[15:8] ? 8'h7d : _GEN_274; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_276 = 8'h14 == io_msg[15:8] ? 8'hfa : _GEN_275; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_277 = 8'h15 == io_msg[15:8] ? 8'h59 : _GEN_276; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_278 = 8'h16 == io_msg[15:8] ? 8'h47 : _GEN_277; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_279 = 8'h17 == io_msg[15:8] ? 8'hf0 : _GEN_278; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_280 = 8'h18 == io_msg[15:8] ? 8'had : _GEN_279; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_281 = 8'h19 == io_msg[15:8] ? 8'hd4 : _GEN_280; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_282 = 8'h1a == io_msg[15:8] ? 8'ha2 : _GEN_281; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_283 = 8'h1b == io_msg[15:8] ? 8'haf : _GEN_282; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_284 = 8'h1c == io_msg[15:8] ? 8'h9c : _GEN_283; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_285 = 8'h1d == io_msg[15:8] ? 8'ha4 : _GEN_284; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_286 = 8'h1e == io_msg[15:8] ? 8'h72 : _GEN_285; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_287 = 8'h1f == io_msg[15:8] ? 8'hc0 : _GEN_286; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_288 = 8'h20 == io_msg[15:8] ? 8'hb7 : _GEN_287; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_289 = 8'h21 == io_msg[15:8] ? 8'hfd : _GEN_288; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_290 = 8'h22 == io_msg[15:8] ? 8'h93 : _GEN_289; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_291 = 8'h23 == io_msg[15:8] ? 8'h26 : _GEN_290; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_292 = 8'h24 == io_msg[15:8] ? 8'h36 : _GEN_291; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_293 = 8'h25 == io_msg[15:8] ? 8'h3f : _GEN_292; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_294 = 8'h26 == io_msg[15:8] ? 8'hf7 : _GEN_293; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_295 = 8'h27 == io_msg[15:8] ? 8'hcc : _GEN_294; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_296 = 8'h28 == io_msg[15:8] ? 8'h34 : _GEN_295; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_297 = 8'h29 == io_msg[15:8] ? 8'ha5 : _GEN_296; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_298 = 8'h2a == io_msg[15:8] ? 8'he5 : _GEN_297; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_299 = 8'h2b == io_msg[15:8] ? 8'hf1 : _GEN_298; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_300 = 8'h2c == io_msg[15:8] ? 8'h71 : _GEN_299; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_301 = 8'h2d == io_msg[15:8] ? 8'hd8 : _GEN_300; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_302 = 8'h2e == io_msg[15:8] ? 8'h31 : _GEN_301; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_303 = 8'h2f == io_msg[15:8] ? 8'h15 : _GEN_302; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_304 = 8'h30 == io_msg[15:8] ? 8'h4 : _GEN_303; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_305 = 8'h31 == io_msg[15:8] ? 8'hc7 : _GEN_304; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_306 = 8'h32 == io_msg[15:8] ? 8'h23 : _GEN_305; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_307 = 8'h33 == io_msg[15:8] ? 8'hc3 : _GEN_306; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_308 = 8'h34 == io_msg[15:8] ? 8'h18 : _GEN_307; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_309 = 8'h35 == io_msg[15:8] ? 8'h96 : _GEN_308; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_310 = 8'h36 == io_msg[15:8] ? 8'h5 : _GEN_309; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_311 = 8'h37 == io_msg[15:8] ? 8'h9a : _GEN_310; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_312 = 8'h38 == io_msg[15:8] ? 8'h7 : _GEN_311; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_313 = 8'h39 == io_msg[15:8] ? 8'h12 : _GEN_312; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_314 = 8'h3a == io_msg[15:8] ? 8'h80 : _GEN_313; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_315 = 8'h3b == io_msg[15:8] ? 8'he2 : _GEN_314; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_316 = 8'h3c == io_msg[15:8] ? 8'heb : _GEN_315; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_317 = 8'h3d == io_msg[15:8] ? 8'h27 : _GEN_316; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_318 = 8'h3e == io_msg[15:8] ? 8'hb2 : _GEN_317; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_319 = 8'h3f == io_msg[15:8] ? 8'h75 : _GEN_318; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_320 = 8'h40 == io_msg[15:8] ? 8'h9 : _GEN_319; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_321 = 8'h41 == io_msg[15:8] ? 8'h83 : _GEN_320; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_322 = 8'h42 == io_msg[15:8] ? 8'h2c : _GEN_321; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_323 = 8'h43 == io_msg[15:8] ? 8'h1a : _GEN_322; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_324 = 8'h44 == io_msg[15:8] ? 8'h1b : _GEN_323; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_325 = 8'h45 == io_msg[15:8] ? 8'h6e : _GEN_324; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_326 = 8'h46 == io_msg[15:8] ? 8'h5a : _GEN_325; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_327 = 8'h47 == io_msg[15:8] ? 8'ha0 : _GEN_326; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_328 = 8'h48 == io_msg[15:8] ? 8'h52 : _GEN_327; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_329 = 8'h49 == io_msg[15:8] ? 8'h3b : _GEN_328; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_330 = 8'h4a == io_msg[15:8] ? 8'hd6 : _GEN_329; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_331 = 8'h4b == io_msg[15:8] ? 8'hb3 : _GEN_330; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_332 = 8'h4c == io_msg[15:8] ? 8'h29 : _GEN_331; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_333 = 8'h4d == io_msg[15:8] ? 8'he3 : _GEN_332; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_334 = 8'h4e == io_msg[15:8] ? 8'h2f : _GEN_333; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_335 = 8'h4f == io_msg[15:8] ? 8'h84 : _GEN_334; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_336 = 8'h50 == io_msg[15:8] ? 8'h53 : _GEN_335; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_337 = 8'h51 == io_msg[15:8] ? 8'hd1 : _GEN_336; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_338 = 8'h52 == io_msg[15:8] ? 8'h0 : _GEN_337; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_339 = 8'h53 == io_msg[15:8] ? 8'hed : _GEN_338; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_340 = 8'h54 == io_msg[15:8] ? 8'h20 : _GEN_339; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_341 = 8'h55 == io_msg[15:8] ? 8'hfc : _GEN_340; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_342 = 8'h56 == io_msg[15:8] ? 8'hb1 : _GEN_341; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_343 = 8'h57 == io_msg[15:8] ? 8'h5b : _GEN_342; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_344 = 8'h58 == io_msg[15:8] ? 8'h6a : _GEN_343; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_345 = 8'h59 == io_msg[15:8] ? 8'hcb : _GEN_344; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_346 = 8'h5a == io_msg[15:8] ? 8'hbe : _GEN_345; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_347 = 8'h5b == io_msg[15:8] ? 8'h39 : _GEN_346; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_348 = 8'h5c == io_msg[15:8] ? 8'h4a : _GEN_347; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_349 = 8'h5d == io_msg[15:8] ? 8'h4c : _GEN_348; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_350 = 8'h5e == io_msg[15:8] ? 8'h58 : _GEN_349; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_351 = 8'h5f == io_msg[15:8] ? 8'hcf : _GEN_350; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_352 = 8'h60 == io_msg[15:8] ? 8'hd0 : _GEN_351; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_353 = 8'h61 == io_msg[15:8] ? 8'hef : _GEN_352; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_354 = 8'h62 == io_msg[15:8] ? 8'haa : _GEN_353; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_355 = 8'h63 == io_msg[15:8] ? 8'hfb : _GEN_354; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_356 = 8'h64 == io_msg[15:8] ? 8'h43 : _GEN_355; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_357 = 8'h65 == io_msg[15:8] ? 8'h4d : _GEN_356; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_358 = 8'h66 == io_msg[15:8] ? 8'h33 : _GEN_357; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_359 = 8'h67 == io_msg[15:8] ? 8'h85 : _GEN_358; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_360 = 8'h68 == io_msg[15:8] ? 8'h45 : _GEN_359; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_361 = 8'h69 == io_msg[15:8] ? 8'hf9 : _GEN_360; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_362 = 8'h6a == io_msg[15:8] ? 8'h2 : _GEN_361; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_363 = 8'h6b == io_msg[15:8] ? 8'h7f : _GEN_362; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_364 = 8'h6c == io_msg[15:8] ? 8'h50 : _GEN_363; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_365 = 8'h6d == io_msg[15:8] ? 8'h3c : _GEN_364; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_366 = 8'h6e == io_msg[15:8] ? 8'h9f : _GEN_365; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_367 = 8'h6f == io_msg[15:8] ? 8'ha8 : _GEN_366; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_368 = 8'h70 == io_msg[15:8] ? 8'h51 : _GEN_367; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_369 = 8'h71 == io_msg[15:8] ? 8'ha3 : _GEN_368; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_370 = 8'h72 == io_msg[15:8] ? 8'h40 : _GEN_369; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_371 = 8'h73 == io_msg[15:8] ? 8'h8f : _GEN_370; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_372 = 8'h74 == io_msg[15:8] ? 8'h92 : _GEN_371; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_373 = 8'h75 == io_msg[15:8] ? 8'h9d : _GEN_372; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_374 = 8'h76 == io_msg[15:8] ? 8'h38 : _GEN_373; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_375 = 8'h77 == io_msg[15:8] ? 8'hf5 : _GEN_374; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_376 = 8'h78 == io_msg[15:8] ? 8'hbc : _GEN_375; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_377 = 8'h79 == io_msg[15:8] ? 8'hb6 : _GEN_376; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_378 = 8'h7a == io_msg[15:8] ? 8'hda : _GEN_377; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_379 = 8'h7b == io_msg[15:8] ? 8'h21 : _GEN_378; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_380 = 8'h7c == io_msg[15:8] ? 8'h10 : _GEN_379; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_381 = 8'h7d == io_msg[15:8] ? 8'hff : _GEN_380; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_382 = 8'h7e == io_msg[15:8] ? 8'hf3 : _GEN_381; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_383 = 8'h7f == io_msg[15:8] ? 8'hd2 : _GEN_382; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_384 = 8'h80 == io_msg[15:8] ? 8'hcd : _GEN_383; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_385 = 8'h81 == io_msg[15:8] ? 8'hc : _GEN_384; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_386 = 8'h82 == io_msg[15:8] ? 8'h13 : _GEN_385; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_387 = 8'h83 == io_msg[15:8] ? 8'hec : _GEN_386; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_388 = 8'h84 == io_msg[15:8] ? 8'h5f : _GEN_387; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_389 = 8'h85 == io_msg[15:8] ? 8'h97 : _GEN_388; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_390 = 8'h86 == io_msg[15:8] ? 8'h44 : _GEN_389; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_391 = 8'h87 == io_msg[15:8] ? 8'h17 : _GEN_390; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_392 = 8'h88 == io_msg[15:8] ? 8'hc4 : _GEN_391; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_393 = 8'h89 == io_msg[15:8] ? 8'ha7 : _GEN_392; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_394 = 8'h8a == io_msg[15:8] ? 8'h7e : _GEN_393; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_395 = 8'h8b == io_msg[15:8] ? 8'h3d : _GEN_394; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_396 = 8'h8c == io_msg[15:8] ? 8'h64 : _GEN_395; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_397 = 8'h8d == io_msg[15:8] ? 8'h5d : _GEN_396; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_398 = 8'h8e == io_msg[15:8] ? 8'h19 : _GEN_397; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_399 = 8'h8f == io_msg[15:8] ? 8'h73 : _GEN_398; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_400 = 8'h90 == io_msg[15:8] ? 8'h60 : _GEN_399; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_401 = 8'h91 == io_msg[15:8] ? 8'h81 : _GEN_400; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_402 = 8'h92 == io_msg[15:8] ? 8'h4f : _GEN_401; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_403 = 8'h93 == io_msg[15:8] ? 8'hdc : _GEN_402; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_404 = 8'h94 == io_msg[15:8] ? 8'h22 : _GEN_403; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_405 = 8'h95 == io_msg[15:8] ? 8'h2a : _GEN_404; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_406 = 8'h96 == io_msg[15:8] ? 8'h90 : _GEN_405; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_407 = 8'h97 == io_msg[15:8] ? 8'h88 : _GEN_406; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_408 = 8'h98 == io_msg[15:8] ? 8'h46 : _GEN_407; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_409 = 8'h99 == io_msg[15:8] ? 8'hee : _GEN_408; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_410 = 8'h9a == io_msg[15:8] ? 8'hb8 : _GEN_409; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_411 = 8'h9b == io_msg[15:8] ? 8'h14 : _GEN_410; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_412 = 8'h9c == io_msg[15:8] ? 8'hde : _GEN_411; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_413 = 8'h9d == io_msg[15:8] ? 8'h5e : _GEN_412; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_414 = 8'h9e == io_msg[15:8] ? 8'hb : _GEN_413; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_415 = 8'h9f == io_msg[15:8] ? 8'hdb : _GEN_414; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_416 = 8'ha0 == io_msg[15:8] ? 8'he0 : _GEN_415; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_417 = 8'ha1 == io_msg[15:8] ? 8'h32 : _GEN_416; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_418 = 8'ha2 == io_msg[15:8] ? 8'h3a : _GEN_417; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_419 = 8'ha3 == io_msg[15:8] ? 8'ha : _GEN_418; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_420 = 8'ha4 == io_msg[15:8] ? 8'h49 : _GEN_419; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_421 = 8'ha5 == io_msg[15:8] ? 8'h6 : _GEN_420; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_422 = 8'ha6 == io_msg[15:8] ? 8'h24 : _GEN_421; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_423 = 8'ha7 == io_msg[15:8] ? 8'h5c : _GEN_422; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_424 = 8'ha8 == io_msg[15:8] ? 8'hc2 : _GEN_423; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_425 = 8'ha9 == io_msg[15:8] ? 8'hd3 : _GEN_424; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_426 = 8'haa == io_msg[15:8] ? 8'hac : _GEN_425; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_427 = 8'hab == io_msg[15:8] ? 8'h62 : _GEN_426; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_428 = 8'hac == io_msg[15:8] ? 8'h91 : _GEN_427; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_429 = 8'had == io_msg[15:8] ? 8'h95 : _GEN_428; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_430 = 8'hae == io_msg[15:8] ? 8'he4 : _GEN_429; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_431 = 8'haf == io_msg[15:8] ? 8'h79 : _GEN_430; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_432 = 8'hb0 == io_msg[15:8] ? 8'he7 : _GEN_431; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_433 = 8'hb1 == io_msg[15:8] ? 8'hc8 : _GEN_432; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_434 = 8'hb2 == io_msg[15:8] ? 8'h37 : _GEN_433; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_435 = 8'hb3 == io_msg[15:8] ? 8'h6d : _GEN_434; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_436 = 8'hb4 == io_msg[15:8] ? 8'h8d : _GEN_435; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_437 = 8'hb5 == io_msg[15:8] ? 8'hd5 : _GEN_436; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_438 = 8'hb6 == io_msg[15:8] ? 8'h4e : _GEN_437; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_439 = 8'hb7 == io_msg[15:8] ? 8'ha9 : _GEN_438; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_440 = 8'hb8 == io_msg[15:8] ? 8'h6c : _GEN_439; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_441 = 8'hb9 == io_msg[15:8] ? 8'h56 : _GEN_440; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_442 = 8'hba == io_msg[15:8] ? 8'hf4 : _GEN_441; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_443 = 8'hbb == io_msg[15:8] ? 8'hea : _GEN_442; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_444 = 8'hbc == io_msg[15:8] ? 8'h65 : _GEN_443; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_445 = 8'hbd == io_msg[15:8] ? 8'h7a : _GEN_444; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_446 = 8'hbe == io_msg[15:8] ? 8'hae : _GEN_445; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_447 = 8'hbf == io_msg[15:8] ? 8'h8 : _GEN_446; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_448 = 8'hc0 == io_msg[15:8] ? 8'hba : _GEN_447; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_449 = 8'hc1 == io_msg[15:8] ? 8'h78 : _GEN_448; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_450 = 8'hc2 == io_msg[15:8] ? 8'h25 : _GEN_449; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_451 = 8'hc3 == io_msg[15:8] ? 8'h2e : _GEN_450; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_452 = 8'hc4 == io_msg[15:8] ? 8'h1c : _GEN_451; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_453 = 8'hc5 == io_msg[15:8] ? 8'ha6 : _GEN_452; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_454 = 8'hc6 == io_msg[15:8] ? 8'hb4 : _GEN_453; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_455 = 8'hc7 == io_msg[15:8] ? 8'hc6 : _GEN_454; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_456 = 8'hc8 == io_msg[15:8] ? 8'he8 : _GEN_455; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_457 = 8'hc9 == io_msg[15:8] ? 8'hdd : _GEN_456; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_458 = 8'hca == io_msg[15:8] ? 8'h74 : _GEN_457; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_459 = 8'hcb == io_msg[15:8] ? 8'h1f : _GEN_458; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_460 = 8'hcc == io_msg[15:8] ? 8'h4b : _GEN_459; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_461 = 8'hcd == io_msg[15:8] ? 8'hbd : _GEN_460; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_462 = 8'hce == io_msg[15:8] ? 8'h8b : _GEN_461; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_463 = 8'hcf == io_msg[15:8] ? 8'h8a : _GEN_462; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_464 = 8'hd0 == io_msg[15:8] ? 8'h70 : _GEN_463; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_465 = 8'hd1 == io_msg[15:8] ? 8'h3e : _GEN_464; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_466 = 8'hd2 == io_msg[15:8] ? 8'hb5 : _GEN_465; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_467 = 8'hd3 == io_msg[15:8] ? 8'h66 : _GEN_466; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_468 = 8'hd4 == io_msg[15:8] ? 8'h48 : _GEN_467; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_469 = 8'hd5 == io_msg[15:8] ? 8'h3 : _GEN_468; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_470 = 8'hd6 == io_msg[15:8] ? 8'hf6 : _GEN_469; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_471 = 8'hd7 == io_msg[15:8] ? 8'he : _GEN_470; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_472 = 8'hd8 == io_msg[15:8] ? 8'h61 : _GEN_471; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_473 = 8'hd9 == io_msg[15:8] ? 8'h35 : _GEN_472; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_474 = 8'hda == io_msg[15:8] ? 8'h57 : _GEN_473; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_475 = 8'hdb == io_msg[15:8] ? 8'hb9 : _GEN_474; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_476 = 8'hdc == io_msg[15:8] ? 8'h86 : _GEN_475; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_477 = 8'hdd == io_msg[15:8] ? 8'hc1 : _GEN_476; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_478 = 8'hde == io_msg[15:8] ? 8'h1d : _GEN_477; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_479 = 8'hdf == io_msg[15:8] ? 8'h9e : _GEN_478; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_480 = 8'he0 == io_msg[15:8] ? 8'he1 : _GEN_479; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_481 = 8'he1 == io_msg[15:8] ? 8'hf8 : _GEN_480; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_482 = 8'he2 == io_msg[15:8] ? 8'h98 : _GEN_481; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_483 = 8'he3 == io_msg[15:8] ? 8'h11 : _GEN_482; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_484 = 8'he4 == io_msg[15:8] ? 8'h69 : _GEN_483; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_485 = 8'he5 == io_msg[15:8] ? 8'hd9 : _GEN_484; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_486 = 8'he6 == io_msg[15:8] ? 8'h8e : _GEN_485; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_487 = 8'he7 == io_msg[15:8] ? 8'h94 : _GEN_486; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_488 = 8'he8 == io_msg[15:8] ? 8'h9b : _GEN_487; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_489 = 8'he9 == io_msg[15:8] ? 8'h1e : _GEN_488; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_490 = 8'hea == io_msg[15:8] ? 8'h87 : _GEN_489; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_491 = 8'heb == io_msg[15:8] ? 8'he9 : _GEN_490; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_492 = 8'hec == io_msg[15:8] ? 8'hce : _GEN_491; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_493 = 8'hed == io_msg[15:8] ? 8'h55 : _GEN_492; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_494 = 8'hee == io_msg[15:8] ? 8'h28 : _GEN_493; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_495 = 8'hef == io_msg[15:8] ? 8'hdf : _GEN_494; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_496 = 8'hf0 == io_msg[15:8] ? 8'h8c : _GEN_495; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_497 = 8'hf1 == io_msg[15:8] ? 8'ha1 : _GEN_496; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_498 = 8'hf2 == io_msg[15:8] ? 8'h89 : _GEN_497; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_499 = 8'hf3 == io_msg[15:8] ? 8'hd : _GEN_498; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_500 = 8'hf4 == io_msg[15:8] ? 8'hbf : _GEN_499; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_501 = 8'hf5 == io_msg[15:8] ? 8'he6 : _GEN_500; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_502 = 8'hf6 == io_msg[15:8] ? 8'h42 : _GEN_501; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_503 = 8'hf7 == io_msg[15:8] ? 8'h68 : _GEN_502; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_504 = 8'hf8 == io_msg[15:8] ? 8'h41 : _GEN_503; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_505 = 8'hf9 == io_msg[15:8] ? 8'h99 : _GEN_504; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_506 = 8'hfa == io_msg[15:8] ? 8'h2d : _GEN_505; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_507 = 8'hfb == io_msg[15:8] ? 8'hf : _GEN_506; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_508 = 8'hfc == io_msg[15:8] ? 8'hb0 : _GEN_507; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_509 = 8'hfd == io_msg[15:8] ? 8'h54 : _GEN_508; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_510 = 8'hfe == io_msg[15:8] ? 8'hbb : _GEN_509; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] sbox_out_1 = 8'hff == io_msg[15:8] ? 8'h16 : _GEN_510; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_513 = 8'h1 == io_msg[23:16] ? 8'h7c : 8'h63; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_514 = 8'h2 == io_msg[23:16] ? 8'h77 : _GEN_513; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_515 = 8'h3 == io_msg[23:16] ? 8'h7b : _GEN_514; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_516 = 8'h4 == io_msg[23:16] ? 8'hf2 : _GEN_515; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_517 = 8'h5 == io_msg[23:16] ? 8'h6b : _GEN_516; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_518 = 8'h6 == io_msg[23:16] ? 8'h6f : _GEN_517; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_519 = 8'h7 == io_msg[23:16] ? 8'hc5 : _GEN_518; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_520 = 8'h8 == io_msg[23:16] ? 8'h30 : _GEN_519; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_521 = 8'h9 == io_msg[23:16] ? 8'h1 : _GEN_520; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_522 = 8'ha == io_msg[23:16] ? 8'h67 : _GEN_521; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_523 = 8'hb == io_msg[23:16] ? 8'h2b : _GEN_522; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_524 = 8'hc == io_msg[23:16] ? 8'hfe : _GEN_523; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_525 = 8'hd == io_msg[23:16] ? 8'hd7 : _GEN_524; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_526 = 8'he == io_msg[23:16] ? 8'hab : _GEN_525; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_527 = 8'hf == io_msg[23:16] ? 8'h76 : _GEN_526; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_528 = 8'h10 == io_msg[23:16] ? 8'hca : _GEN_527; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_529 = 8'h11 == io_msg[23:16] ? 8'h82 : _GEN_528; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_530 = 8'h12 == io_msg[23:16] ? 8'hc9 : _GEN_529; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_531 = 8'h13 == io_msg[23:16] ? 8'h7d : _GEN_530; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_532 = 8'h14 == io_msg[23:16] ? 8'hfa : _GEN_531; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_533 = 8'h15 == io_msg[23:16] ? 8'h59 : _GEN_532; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_534 = 8'h16 == io_msg[23:16] ? 8'h47 : _GEN_533; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_535 = 8'h17 == io_msg[23:16] ? 8'hf0 : _GEN_534; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_536 = 8'h18 == io_msg[23:16] ? 8'had : _GEN_535; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_537 = 8'h19 == io_msg[23:16] ? 8'hd4 : _GEN_536; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_538 = 8'h1a == io_msg[23:16] ? 8'ha2 : _GEN_537; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_539 = 8'h1b == io_msg[23:16] ? 8'haf : _GEN_538; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_540 = 8'h1c == io_msg[23:16] ? 8'h9c : _GEN_539; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_541 = 8'h1d == io_msg[23:16] ? 8'ha4 : _GEN_540; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_542 = 8'h1e == io_msg[23:16] ? 8'h72 : _GEN_541; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_543 = 8'h1f == io_msg[23:16] ? 8'hc0 : _GEN_542; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_544 = 8'h20 == io_msg[23:16] ? 8'hb7 : _GEN_543; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_545 = 8'h21 == io_msg[23:16] ? 8'hfd : _GEN_544; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_546 = 8'h22 == io_msg[23:16] ? 8'h93 : _GEN_545; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_547 = 8'h23 == io_msg[23:16] ? 8'h26 : _GEN_546; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_548 = 8'h24 == io_msg[23:16] ? 8'h36 : _GEN_547; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_549 = 8'h25 == io_msg[23:16] ? 8'h3f : _GEN_548; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_550 = 8'h26 == io_msg[23:16] ? 8'hf7 : _GEN_549; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_551 = 8'h27 == io_msg[23:16] ? 8'hcc : _GEN_550; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_552 = 8'h28 == io_msg[23:16] ? 8'h34 : _GEN_551; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_553 = 8'h29 == io_msg[23:16] ? 8'ha5 : _GEN_552; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_554 = 8'h2a == io_msg[23:16] ? 8'he5 : _GEN_553; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_555 = 8'h2b == io_msg[23:16] ? 8'hf1 : _GEN_554; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_556 = 8'h2c == io_msg[23:16] ? 8'h71 : _GEN_555; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_557 = 8'h2d == io_msg[23:16] ? 8'hd8 : _GEN_556; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_558 = 8'h2e == io_msg[23:16] ? 8'h31 : _GEN_557; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_559 = 8'h2f == io_msg[23:16] ? 8'h15 : _GEN_558; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_560 = 8'h30 == io_msg[23:16] ? 8'h4 : _GEN_559; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_561 = 8'h31 == io_msg[23:16] ? 8'hc7 : _GEN_560; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_562 = 8'h32 == io_msg[23:16] ? 8'h23 : _GEN_561; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_563 = 8'h33 == io_msg[23:16] ? 8'hc3 : _GEN_562; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_564 = 8'h34 == io_msg[23:16] ? 8'h18 : _GEN_563; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_565 = 8'h35 == io_msg[23:16] ? 8'h96 : _GEN_564; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_566 = 8'h36 == io_msg[23:16] ? 8'h5 : _GEN_565; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_567 = 8'h37 == io_msg[23:16] ? 8'h9a : _GEN_566; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_568 = 8'h38 == io_msg[23:16] ? 8'h7 : _GEN_567; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_569 = 8'h39 == io_msg[23:16] ? 8'h12 : _GEN_568; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_570 = 8'h3a == io_msg[23:16] ? 8'h80 : _GEN_569; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_571 = 8'h3b == io_msg[23:16] ? 8'he2 : _GEN_570; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_572 = 8'h3c == io_msg[23:16] ? 8'heb : _GEN_571; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_573 = 8'h3d == io_msg[23:16] ? 8'h27 : _GEN_572; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_574 = 8'h3e == io_msg[23:16] ? 8'hb2 : _GEN_573; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_575 = 8'h3f == io_msg[23:16] ? 8'h75 : _GEN_574; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_576 = 8'h40 == io_msg[23:16] ? 8'h9 : _GEN_575; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_577 = 8'h41 == io_msg[23:16] ? 8'h83 : _GEN_576; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_578 = 8'h42 == io_msg[23:16] ? 8'h2c : _GEN_577; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_579 = 8'h43 == io_msg[23:16] ? 8'h1a : _GEN_578; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_580 = 8'h44 == io_msg[23:16] ? 8'h1b : _GEN_579; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_581 = 8'h45 == io_msg[23:16] ? 8'h6e : _GEN_580; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_582 = 8'h46 == io_msg[23:16] ? 8'h5a : _GEN_581; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_583 = 8'h47 == io_msg[23:16] ? 8'ha0 : _GEN_582; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_584 = 8'h48 == io_msg[23:16] ? 8'h52 : _GEN_583; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_585 = 8'h49 == io_msg[23:16] ? 8'h3b : _GEN_584; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_586 = 8'h4a == io_msg[23:16] ? 8'hd6 : _GEN_585; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_587 = 8'h4b == io_msg[23:16] ? 8'hb3 : _GEN_586; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_588 = 8'h4c == io_msg[23:16] ? 8'h29 : _GEN_587; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_589 = 8'h4d == io_msg[23:16] ? 8'he3 : _GEN_588; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_590 = 8'h4e == io_msg[23:16] ? 8'h2f : _GEN_589; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_591 = 8'h4f == io_msg[23:16] ? 8'h84 : _GEN_590; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_592 = 8'h50 == io_msg[23:16] ? 8'h53 : _GEN_591; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_593 = 8'h51 == io_msg[23:16] ? 8'hd1 : _GEN_592; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_594 = 8'h52 == io_msg[23:16] ? 8'h0 : _GEN_593; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_595 = 8'h53 == io_msg[23:16] ? 8'hed : _GEN_594; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_596 = 8'h54 == io_msg[23:16] ? 8'h20 : _GEN_595; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_597 = 8'h55 == io_msg[23:16] ? 8'hfc : _GEN_596; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_598 = 8'h56 == io_msg[23:16] ? 8'hb1 : _GEN_597; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_599 = 8'h57 == io_msg[23:16] ? 8'h5b : _GEN_598; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_600 = 8'h58 == io_msg[23:16] ? 8'h6a : _GEN_599; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_601 = 8'h59 == io_msg[23:16] ? 8'hcb : _GEN_600; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_602 = 8'h5a == io_msg[23:16] ? 8'hbe : _GEN_601; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_603 = 8'h5b == io_msg[23:16] ? 8'h39 : _GEN_602; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_604 = 8'h5c == io_msg[23:16] ? 8'h4a : _GEN_603; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_605 = 8'h5d == io_msg[23:16] ? 8'h4c : _GEN_604; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_606 = 8'h5e == io_msg[23:16] ? 8'h58 : _GEN_605; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_607 = 8'h5f == io_msg[23:16] ? 8'hcf : _GEN_606; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_608 = 8'h60 == io_msg[23:16] ? 8'hd0 : _GEN_607; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_609 = 8'h61 == io_msg[23:16] ? 8'hef : _GEN_608; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_610 = 8'h62 == io_msg[23:16] ? 8'haa : _GEN_609; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_611 = 8'h63 == io_msg[23:16] ? 8'hfb : _GEN_610; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_612 = 8'h64 == io_msg[23:16] ? 8'h43 : _GEN_611; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_613 = 8'h65 == io_msg[23:16] ? 8'h4d : _GEN_612; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_614 = 8'h66 == io_msg[23:16] ? 8'h33 : _GEN_613; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_615 = 8'h67 == io_msg[23:16] ? 8'h85 : _GEN_614; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_616 = 8'h68 == io_msg[23:16] ? 8'h45 : _GEN_615; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_617 = 8'h69 == io_msg[23:16] ? 8'hf9 : _GEN_616; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_618 = 8'h6a == io_msg[23:16] ? 8'h2 : _GEN_617; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_619 = 8'h6b == io_msg[23:16] ? 8'h7f : _GEN_618; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_620 = 8'h6c == io_msg[23:16] ? 8'h50 : _GEN_619; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_621 = 8'h6d == io_msg[23:16] ? 8'h3c : _GEN_620; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_622 = 8'h6e == io_msg[23:16] ? 8'h9f : _GEN_621; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_623 = 8'h6f == io_msg[23:16] ? 8'ha8 : _GEN_622; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_624 = 8'h70 == io_msg[23:16] ? 8'h51 : _GEN_623; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_625 = 8'h71 == io_msg[23:16] ? 8'ha3 : _GEN_624; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_626 = 8'h72 == io_msg[23:16] ? 8'h40 : _GEN_625; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_627 = 8'h73 == io_msg[23:16] ? 8'h8f : _GEN_626; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_628 = 8'h74 == io_msg[23:16] ? 8'h92 : _GEN_627; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_629 = 8'h75 == io_msg[23:16] ? 8'h9d : _GEN_628; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_630 = 8'h76 == io_msg[23:16] ? 8'h38 : _GEN_629; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_631 = 8'h77 == io_msg[23:16] ? 8'hf5 : _GEN_630; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_632 = 8'h78 == io_msg[23:16] ? 8'hbc : _GEN_631; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_633 = 8'h79 == io_msg[23:16] ? 8'hb6 : _GEN_632; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_634 = 8'h7a == io_msg[23:16] ? 8'hda : _GEN_633; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_635 = 8'h7b == io_msg[23:16] ? 8'h21 : _GEN_634; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_636 = 8'h7c == io_msg[23:16] ? 8'h10 : _GEN_635; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_637 = 8'h7d == io_msg[23:16] ? 8'hff : _GEN_636; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_638 = 8'h7e == io_msg[23:16] ? 8'hf3 : _GEN_637; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_639 = 8'h7f == io_msg[23:16] ? 8'hd2 : _GEN_638; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_640 = 8'h80 == io_msg[23:16] ? 8'hcd : _GEN_639; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_641 = 8'h81 == io_msg[23:16] ? 8'hc : _GEN_640; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_642 = 8'h82 == io_msg[23:16] ? 8'h13 : _GEN_641; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_643 = 8'h83 == io_msg[23:16] ? 8'hec : _GEN_642; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_644 = 8'h84 == io_msg[23:16] ? 8'h5f : _GEN_643; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_645 = 8'h85 == io_msg[23:16] ? 8'h97 : _GEN_644; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_646 = 8'h86 == io_msg[23:16] ? 8'h44 : _GEN_645; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_647 = 8'h87 == io_msg[23:16] ? 8'h17 : _GEN_646; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_648 = 8'h88 == io_msg[23:16] ? 8'hc4 : _GEN_647; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_649 = 8'h89 == io_msg[23:16] ? 8'ha7 : _GEN_648; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_650 = 8'h8a == io_msg[23:16] ? 8'h7e : _GEN_649; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_651 = 8'h8b == io_msg[23:16] ? 8'h3d : _GEN_650; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_652 = 8'h8c == io_msg[23:16] ? 8'h64 : _GEN_651; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_653 = 8'h8d == io_msg[23:16] ? 8'h5d : _GEN_652; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_654 = 8'h8e == io_msg[23:16] ? 8'h19 : _GEN_653; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_655 = 8'h8f == io_msg[23:16] ? 8'h73 : _GEN_654; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_656 = 8'h90 == io_msg[23:16] ? 8'h60 : _GEN_655; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_657 = 8'h91 == io_msg[23:16] ? 8'h81 : _GEN_656; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_658 = 8'h92 == io_msg[23:16] ? 8'h4f : _GEN_657; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_659 = 8'h93 == io_msg[23:16] ? 8'hdc : _GEN_658; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_660 = 8'h94 == io_msg[23:16] ? 8'h22 : _GEN_659; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_661 = 8'h95 == io_msg[23:16] ? 8'h2a : _GEN_660; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_662 = 8'h96 == io_msg[23:16] ? 8'h90 : _GEN_661; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_663 = 8'h97 == io_msg[23:16] ? 8'h88 : _GEN_662; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_664 = 8'h98 == io_msg[23:16] ? 8'h46 : _GEN_663; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_665 = 8'h99 == io_msg[23:16] ? 8'hee : _GEN_664; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_666 = 8'h9a == io_msg[23:16] ? 8'hb8 : _GEN_665; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_667 = 8'h9b == io_msg[23:16] ? 8'h14 : _GEN_666; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_668 = 8'h9c == io_msg[23:16] ? 8'hde : _GEN_667; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_669 = 8'h9d == io_msg[23:16] ? 8'h5e : _GEN_668; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_670 = 8'h9e == io_msg[23:16] ? 8'hb : _GEN_669; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_671 = 8'h9f == io_msg[23:16] ? 8'hdb : _GEN_670; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_672 = 8'ha0 == io_msg[23:16] ? 8'he0 : _GEN_671; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_673 = 8'ha1 == io_msg[23:16] ? 8'h32 : _GEN_672; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_674 = 8'ha2 == io_msg[23:16] ? 8'h3a : _GEN_673; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_675 = 8'ha3 == io_msg[23:16] ? 8'ha : _GEN_674; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_676 = 8'ha4 == io_msg[23:16] ? 8'h49 : _GEN_675; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_677 = 8'ha5 == io_msg[23:16] ? 8'h6 : _GEN_676; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_678 = 8'ha6 == io_msg[23:16] ? 8'h24 : _GEN_677; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_679 = 8'ha7 == io_msg[23:16] ? 8'h5c : _GEN_678; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_680 = 8'ha8 == io_msg[23:16] ? 8'hc2 : _GEN_679; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_681 = 8'ha9 == io_msg[23:16] ? 8'hd3 : _GEN_680; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_682 = 8'haa == io_msg[23:16] ? 8'hac : _GEN_681; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_683 = 8'hab == io_msg[23:16] ? 8'h62 : _GEN_682; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_684 = 8'hac == io_msg[23:16] ? 8'h91 : _GEN_683; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_685 = 8'had == io_msg[23:16] ? 8'h95 : _GEN_684; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_686 = 8'hae == io_msg[23:16] ? 8'he4 : _GEN_685; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_687 = 8'haf == io_msg[23:16] ? 8'h79 : _GEN_686; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_688 = 8'hb0 == io_msg[23:16] ? 8'he7 : _GEN_687; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_689 = 8'hb1 == io_msg[23:16] ? 8'hc8 : _GEN_688; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_690 = 8'hb2 == io_msg[23:16] ? 8'h37 : _GEN_689; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_691 = 8'hb3 == io_msg[23:16] ? 8'h6d : _GEN_690; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_692 = 8'hb4 == io_msg[23:16] ? 8'h8d : _GEN_691; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_693 = 8'hb5 == io_msg[23:16] ? 8'hd5 : _GEN_692; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_694 = 8'hb6 == io_msg[23:16] ? 8'h4e : _GEN_693; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_695 = 8'hb7 == io_msg[23:16] ? 8'ha9 : _GEN_694; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_696 = 8'hb8 == io_msg[23:16] ? 8'h6c : _GEN_695; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_697 = 8'hb9 == io_msg[23:16] ? 8'h56 : _GEN_696; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_698 = 8'hba == io_msg[23:16] ? 8'hf4 : _GEN_697; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_699 = 8'hbb == io_msg[23:16] ? 8'hea : _GEN_698; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_700 = 8'hbc == io_msg[23:16] ? 8'h65 : _GEN_699; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_701 = 8'hbd == io_msg[23:16] ? 8'h7a : _GEN_700; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_702 = 8'hbe == io_msg[23:16] ? 8'hae : _GEN_701; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_703 = 8'hbf == io_msg[23:16] ? 8'h8 : _GEN_702; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_704 = 8'hc0 == io_msg[23:16] ? 8'hba : _GEN_703; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_705 = 8'hc1 == io_msg[23:16] ? 8'h78 : _GEN_704; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_706 = 8'hc2 == io_msg[23:16] ? 8'h25 : _GEN_705; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_707 = 8'hc3 == io_msg[23:16] ? 8'h2e : _GEN_706; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_708 = 8'hc4 == io_msg[23:16] ? 8'h1c : _GEN_707; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_709 = 8'hc5 == io_msg[23:16] ? 8'ha6 : _GEN_708; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_710 = 8'hc6 == io_msg[23:16] ? 8'hb4 : _GEN_709; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_711 = 8'hc7 == io_msg[23:16] ? 8'hc6 : _GEN_710; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_712 = 8'hc8 == io_msg[23:16] ? 8'he8 : _GEN_711; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_713 = 8'hc9 == io_msg[23:16] ? 8'hdd : _GEN_712; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_714 = 8'hca == io_msg[23:16] ? 8'h74 : _GEN_713; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_715 = 8'hcb == io_msg[23:16] ? 8'h1f : _GEN_714; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_716 = 8'hcc == io_msg[23:16] ? 8'h4b : _GEN_715; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_717 = 8'hcd == io_msg[23:16] ? 8'hbd : _GEN_716; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_718 = 8'hce == io_msg[23:16] ? 8'h8b : _GEN_717; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_719 = 8'hcf == io_msg[23:16] ? 8'h8a : _GEN_718; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_720 = 8'hd0 == io_msg[23:16] ? 8'h70 : _GEN_719; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_721 = 8'hd1 == io_msg[23:16] ? 8'h3e : _GEN_720; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_722 = 8'hd2 == io_msg[23:16] ? 8'hb5 : _GEN_721; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_723 = 8'hd3 == io_msg[23:16] ? 8'h66 : _GEN_722; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_724 = 8'hd4 == io_msg[23:16] ? 8'h48 : _GEN_723; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_725 = 8'hd5 == io_msg[23:16] ? 8'h3 : _GEN_724; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_726 = 8'hd6 == io_msg[23:16] ? 8'hf6 : _GEN_725; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_727 = 8'hd7 == io_msg[23:16] ? 8'he : _GEN_726; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_728 = 8'hd8 == io_msg[23:16] ? 8'h61 : _GEN_727; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_729 = 8'hd9 == io_msg[23:16] ? 8'h35 : _GEN_728; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_730 = 8'hda == io_msg[23:16] ? 8'h57 : _GEN_729; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_731 = 8'hdb == io_msg[23:16] ? 8'hb9 : _GEN_730; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_732 = 8'hdc == io_msg[23:16] ? 8'h86 : _GEN_731; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_733 = 8'hdd == io_msg[23:16] ? 8'hc1 : _GEN_732; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_734 = 8'hde == io_msg[23:16] ? 8'h1d : _GEN_733; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_735 = 8'hdf == io_msg[23:16] ? 8'h9e : _GEN_734; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_736 = 8'he0 == io_msg[23:16] ? 8'he1 : _GEN_735; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_737 = 8'he1 == io_msg[23:16] ? 8'hf8 : _GEN_736; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_738 = 8'he2 == io_msg[23:16] ? 8'h98 : _GEN_737; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_739 = 8'he3 == io_msg[23:16] ? 8'h11 : _GEN_738; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_740 = 8'he4 == io_msg[23:16] ? 8'h69 : _GEN_739; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_741 = 8'he5 == io_msg[23:16] ? 8'hd9 : _GEN_740; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_742 = 8'he6 == io_msg[23:16] ? 8'h8e : _GEN_741; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_743 = 8'he7 == io_msg[23:16] ? 8'h94 : _GEN_742; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_744 = 8'he8 == io_msg[23:16] ? 8'h9b : _GEN_743; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_745 = 8'he9 == io_msg[23:16] ? 8'h1e : _GEN_744; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_746 = 8'hea == io_msg[23:16] ? 8'h87 : _GEN_745; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_747 = 8'heb == io_msg[23:16] ? 8'he9 : _GEN_746; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_748 = 8'hec == io_msg[23:16] ? 8'hce : _GEN_747; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_749 = 8'hed == io_msg[23:16] ? 8'h55 : _GEN_748; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_750 = 8'hee == io_msg[23:16] ? 8'h28 : _GEN_749; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_751 = 8'hef == io_msg[23:16] ? 8'hdf : _GEN_750; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_752 = 8'hf0 == io_msg[23:16] ? 8'h8c : _GEN_751; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_753 = 8'hf1 == io_msg[23:16] ? 8'ha1 : _GEN_752; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_754 = 8'hf2 == io_msg[23:16] ? 8'h89 : _GEN_753; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_755 = 8'hf3 == io_msg[23:16] ? 8'hd : _GEN_754; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_756 = 8'hf4 == io_msg[23:16] ? 8'hbf : _GEN_755; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_757 = 8'hf5 == io_msg[23:16] ? 8'he6 : _GEN_756; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_758 = 8'hf6 == io_msg[23:16] ? 8'h42 : _GEN_757; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_759 = 8'hf7 == io_msg[23:16] ? 8'h68 : _GEN_758; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_760 = 8'hf8 == io_msg[23:16] ? 8'h41 : _GEN_759; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_761 = 8'hf9 == io_msg[23:16] ? 8'h99 : _GEN_760; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_762 = 8'hfa == io_msg[23:16] ? 8'h2d : _GEN_761; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_763 = 8'hfb == io_msg[23:16] ? 8'hf : _GEN_762; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_764 = 8'hfc == io_msg[23:16] ? 8'hb0 : _GEN_763; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_765 = 8'hfd == io_msg[23:16] ? 8'h54 : _GEN_764; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_766 = 8'hfe == io_msg[23:16] ? 8'hbb : _GEN_765; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] sbox_out_2 = 8'hff == io_msg[23:16] ? 8'h16 : _GEN_766; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_769 = 8'h1 == io_msg[31:24] ? 8'h7c : 8'h63; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_770 = 8'h2 == io_msg[31:24] ? 8'h77 : _GEN_769; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_771 = 8'h3 == io_msg[31:24] ? 8'h7b : _GEN_770; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_772 = 8'h4 == io_msg[31:24] ? 8'hf2 : _GEN_771; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_773 = 8'h5 == io_msg[31:24] ? 8'h6b : _GEN_772; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_774 = 8'h6 == io_msg[31:24] ? 8'h6f : _GEN_773; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_775 = 8'h7 == io_msg[31:24] ? 8'hc5 : _GEN_774; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_776 = 8'h8 == io_msg[31:24] ? 8'h30 : _GEN_775; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_777 = 8'h9 == io_msg[31:24] ? 8'h1 : _GEN_776; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_778 = 8'ha == io_msg[31:24] ? 8'h67 : _GEN_777; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_779 = 8'hb == io_msg[31:24] ? 8'h2b : _GEN_778; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_780 = 8'hc == io_msg[31:24] ? 8'hfe : _GEN_779; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_781 = 8'hd == io_msg[31:24] ? 8'hd7 : _GEN_780; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_782 = 8'he == io_msg[31:24] ? 8'hab : _GEN_781; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_783 = 8'hf == io_msg[31:24] ? 8'h76 : _GEN_782; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_784 = 8'h10 == io_msg[31:24] ? 8'hca : _GEN_783; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_785 = 8'h11 == io_msg[31:24] ? 8'h82 : _GEN_784; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_786 = 8'h12 == io_msg[31:24] ? 8'hc9 : _GEN_785; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_787 = 8'h13 == io_msg[31:24] ? 8'h7d : _GEN_786; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_788 = 8'h14 == io_msg[31:24] ? 8'hfa : _GEN_787; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_789 = 8'h15 == io_msg[31:24] ? 8'h59 : _GEN_788; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_790 = 8'h16 == io_msg[31:24] ? 8'h47 : _GEN_789; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_791 = 8'h17 == io_msg[31:24] ? 8'hf0 : _GEN_790; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_792 = 8'h18 == io_msg[31:24] ? 8'had : _GEN_791; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_793 = 8'h19 == io_msg[31:24] ? 8'hd4 : _GEN_792; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_794 = 8'h1a == io_msg[31:24] ? 8'ha2 : _GEN_793; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_795 = 8'h1b == io_msg[31:24] ? 8'haf : _GEN_794; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_796 = 8'h1c == io_msg[31:24] ? 8'h9c : _GEN_795; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_797 = 8'h1d == io_msg[31:24] ? 8'ha4 : _GEN_796; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_798 = 8'h1e == io_msg[31:24] ? 8'h72 : _GEN_797; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_799 = 8'h1f == io_msg[31:24] ? 8'hc0 : _GEN_798; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_800 = 8'h20 == io_msg[31:24] ? 8'hb7 : _GEN_799; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_801 = 8'h21 == io_msg[31:24] ? 8'hfd : _GEN_800; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_802 = 8'h22 == io_msg[31:24] ? 8'h93 : _GEN_801; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_803 = 8'h23 == io_msg[31:24] ? 8'h26 : _GEN_802; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_804 = 8'h24 == io_msg[31:24] ? 8'h36 : _GEN_803; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_805 = 8'h25 == io_msg[31:24] ? 8'h3f : _GEN_804; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_806 = 8'h26 == io_msg[31:24] ? 8'hf7 : _GEN_805; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_807 = 8'h27 == io_msg[31:24] ? 8'hcc : _GEN_806; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_808 = 8'h28 == io_msg[31:24] ? 8'h34 : _GEN_807; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_809 = 8'h29 == io_msg[31:24] ? 8'ha5 : _GEN_808; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_810 = 8'h2a == io_msg[31:24] ? 8'he5 : _GEN_809; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_811 = 8'h2b == io_msg[31:24] ? 8'hf1 : _GEN_810; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_812 = 8'h2c == io_msg[31:24] ? 8'h71 : _GEN_811; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_813 = 8'h2d == io_msg[31:24] ? 8'hd8 : _GEN_812; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_814 = 8'h2e == io_msg[31:24] ? 8'h31 : _GEN_813; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_815 = 8'h2f == io_msg[31:24] ? 8'h15 : _GEN_814; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_816 = 8'h30 == io_msg[31:24] ? 8'h4 : _GEN_815; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_817 = 8'h31 == io_msg[31:24] ? 8'hc7 : _GEN_816; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_818 = 8'h32 == io_msg[31:24] ? 8'h23 : _GEN_817; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_819 = 8'h33 == io_msg[31:24] ? 8'hc3 : _GEN_818; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_820 = 8'h34 == io_msg[31:24] ? 8'h18 : _GEN_819; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_821 = 8'h35 == io_msg[31:24] ? 8'h96 : _GEN_820; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_822 = 8'h36 == io_msg[31:24] ? 8'h5 : _GEN_821; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_823 = 8'h37 == io_msg[31:24] ? 8'h9a : _GEN_822; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_824 = 8'h38 == io_msg[31:24] ? 8'h7 : _GEN_823; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_825 = 8'h39 == io_msg[31:24] ? 8'h12 : _GEN_824; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_826 = 8'h3a == io_msg[31:24] ? 8'h80 : _GEN_825; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_827 = 8'h3b == io_msg[31:24] ? 8'he2 : _GEN_826; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_828 = 8'h3c == io_msg[31:24] ? 8'heb : _GEN_827; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_829 = 8'h3d == io_msg[31:24] ? 8'h27 : _GEN_828; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_830 = 8'h3e == io_msg[31:24] ? 8'hb2 : _GEN_829; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_831 = 8'h3f == io_msg[31:24] ? 8'h75 : _GEN_830; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_832 = 8'h40 == io_msg[31:24] ? 8'h9 : _GEN_831; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_833 = 8'h41 == io_msg[31:24] ? 8'h83 : _GEN_832; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_834 = 8'h42 == io_msg[31:24] ? 8'h2c : _GEN_833; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_835 = 8'h43 == io_msg[31:24] ? 8'h1a : _GEN_834; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_836 = 8'h44 == io_msg[31:24] ? 8'h1b : _GEN_835; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_837 = 8'h45 == io_msg[31:24] ? 8'h6e : _GEN_836; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_838 = 8'h46 == io_msg[31:24] ? 8'h5a : _GEN_837; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_839 = 8'h47 == io_msg[31:24] ? 8'ha0 : _GEN_838; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_840 = 8'h48 == io_msg[31:24] ? 8'h52 : _GEN_839; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_841 = 8'h49 == io_msg[31:24] ? 8'h3b : _GEN_840; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_842 = 8'h4a == io_msg[31:24] ? 8'hd6 : _GEN_841; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_843 = 8'h4b == io_msg[31:24] ? 8'hb3 : _GEN_842; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_844 = 8'h4c == io_msg[31:24] ? 8'h29 : _GEN_843; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_845 = 8'h4d == io_msg[31:24] ? 8'he3 : _GEN_844; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_846 = 8'h4e == io_msg[31:24] ? 8'h2f : _GEN_845; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_847 = 8'h4f == io_msg[31:24] ? 8'h84 : _GEN_846; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_848 = 8'h50 == io_msg[31:24] ? 8'h53 : _GEN_847; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_849 = 8'h51 == io_msg[31:24] ? 8'hd1 : _GEN_848; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_850 = 8'h52 == io_msg[31:24] ? 8'h0 : _GEN_849; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_851 = 8'h53 == io_msg[31:24] ? 8'hed : _GEN_850; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_852 = 8'h54 == io_msg[31:24] ? 8'h20 : _GEN_851; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_853 = 8'h55 == io_msg[31:24] ? 8'hfc : _GEN_852; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_854 = 8'h56 == io_msg[31:24] ? 8'hb1 : _GEN_853; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_855 = 8'h57 == io_msg[31:24] ? 8'h5b : _GEN_854; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_856 = 8'h58 == io_msg[31:24] ? 8'h6a : _GEN_855; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_857 = 8'h59 == io_msg[31:24] ? 8'hcb : _GEN_856; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_858 = 8'h5a == io_msg[31:24] ? 8'hbe : _GEN_857; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_859 = 8'h5b == io_msg[31:24] ? 8'h39 : _GEN_858; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_860 = 8'h5c == io_msg[31:24] ? 8'h4a : _GEN_859; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_861 = 8'h5d == io_msg[31:24] ? 8'h4c : _GEN_860; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_862 = 8'h5e == io_msg[31:24] ? 8'h58 : _GEN_861; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_863 = 8'h5f == io_msg[31:24] ? 8'hcf : _GEN_862; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_864 = 8'h60 == io_msg[31:24] ? 8'hd0 : _GEN_863; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_865 = 8'h61 == io_msg[31:24] ? 8'hef : _GEN_864; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_866 = 8'h62 == io_msg[31:24] ? 8'haa : _GEN_865; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_867 = 8'h63 == io_msg[31:24] ? 8'hfb : _GEN_866; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_868 = 8'h64 == io_msg[31:24] ? 8'h43 : _GEN_867; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_869 = 8'h65 == io_msg[31:24] ? 8'h4d : _GEN_868; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_870 = 8'h66 == io_msg[31:24] ? 8'h33 : _GEN_869; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_871 = 8'h67 == io_msg[31:24] ? 8'h85 : _GEN_870; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_872 = 8'h68 == io_msg[31:24] ? 8'h45 : _GEN_871; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_873 = 8'h69 == io_msg[31:24] ? 8'hf9 : _GEN_872; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_874 = 8'h6a == io_msg[31:24] ? 8'h2 : _GEN_873; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_875 = 8'h6b == io_msg[31:24] ? 8'h7f : _GEN_874; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_876 = 8'h6c == io_msg[31:24] ? 8'h50 : _GEN_875; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_877 = 8'h6d == io_msg[31:24] ? 8'h3c : _GEN_876; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_878 = 8'h6e == io_msg[31:24] ? 8'h9f : _GEN_877; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_879 = 8'h6f == io_msg[31:24] ? 8'ha8 : _GEN_878; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_880 = 8'h70 == io_msg[31:24] ? 8'h51 : _GEN_879; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_881 = 8'h71 == io_msg[31:24] ? 8'ha3 : _GEN_880; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_882 = 8'h72 == io_msg[31:24] ? 8'h40 : _GEN_881; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_883 = 8'h73 == io_msg[31:24] ? 8'h8f : _GEN_882; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_884 = 8'h74 == io_msg[31:24] ? 8'h92 : _GEN_883; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_885 = 8'h75 == io_msg[31:24] ? 8'h9d : _GEN_884; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_886 = 8'h76 == io_msg[31:24] ? 8'h38 : _GEN_885; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_887 = 8'h77 == io_msg[31:24] ? 8'hf5 : _GEN_886; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_888 = 8'h78 == io_msg[31:24] ? 8'hbc : _GEN_887; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_889 = 8'h79 == io_msg[31:24] ? 8'hb6 : _GEN_888; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_890 = 8'h7a == io_msg[31:24] ? 8'hda : _GEN_889; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_891 = 8'h7b == io_msg[31:24] ? 8'h21 : _GEN_890; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_892 = 8'h7c == io_msg[31:24] ? 8'h10 : _GEN_891; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_893 = 8'h7d == io_msg[31:24] ? 8'hff : _GEN_892; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_894 = 8'h7e == io_msg[31:24] ? 8'hf3 : _GEN_893; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_895 = 8'h7f == io_msg[31:24] ? 8'hd2 : _GEN_894; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_896 = 8'h80 == io_msg[31:24] ? 8'hcd : _GEN_895; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_897 = 8'h81 == io_msg[31:24] ? 8'hc : _GEN_896; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_898 = 8'h82 == io_msg[31:24] ? 8'h13 : _GEN_897; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_899 = 8'h83 == io_msg[31:24] ? 8'hec : _GEN_898; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_900 = 8'h84 == io_msg[31:24] ? 8'h5f : _GEN_899; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_901 = 8'h85 == io_msg[31:24] ? 8'h97 : _GEN_900; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_902 = 8'h86 == io_msg[31:24] ? 8'h44 : _GEN_901; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_903 = 8'h87 == io_msg[31:24] ? 8'h17 : _GEN_902; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_904 = 8'h88 == io_msg[31:24] ? 8'hc4 : _GEN_903; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_905 = 8'h89 == io_msg[31:24] ? 8'ha7 : _GEN_904; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_906 = 8'h8a == io_msg[31:24] ? 8'h7e : _GEN_905; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_907 = 8'h8b == io_msg[31:24] ? 8'h3d : _GEN_906; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_908 = 8'h8c == io_msg[31:24] ? 8'h64 : _GEN_907; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_909 = 8'h8d == io_msg[31:24] ? 8'h5d : _GEN_908; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_910 = 8'h8e == io_msg[31:24] ? 8'h19 : _GEN_909; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_911 = 8'h8f == io_msg[31:24] ? 8'h73 : _GEN_910; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_912 = 8'h90 == io_msg[31:24] ? 8'h60 : _GEN_911; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_913 = 8'h91 == io_msg[31:24] ? 8'h81 : _GEN_912; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_914 = 8'h92 == io_msg[31:24] ? 8'h4f : _GEN_913; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_915 = 8'h93 == io_msg[31:24] ? 8'hdc : _GEN_914; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_916 = 8'h94 == io_msg[31:24] ? 8'h22 : _GEN_915; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_917 = 8'h95 == io_msg[31:24] ? 8'h2a : _GEN_916; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_918 = 8'h96 == io_msg[31:24] ? 8'h90 : _GEN_917; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_919 = 8'h97 == io_msg[31:24] ? 8'h88 : _GEN_918; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_920 = 8'h98 == io_msg[31:24] ? 8'h46 : _GEN_919; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_921 = 8'h99 == io_msg[31:24] ? 8'hee : _GEN_920; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_922 = 8'h9a == io_msg[31:24] ? 8'hb8 : _GEN_921; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_923 = 8'h9b == io_msg[31:24] ? 8'h14 : _GEN_922; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_924 = 8'h9c == io_msg[31:24] ? 8'hde : _GEN_923; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_925 = 8'h9d == io_msg[31:24] ? 8'h5e : _GEN_924; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_926 = 8'h9e == io_msg[31:24] ? 8'hb : _GEN_925; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_927 = 8'h9f == io_msg[31:24] ? 8'hdb : _GEN_926; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_928 = 8'ha0 == io_msg[31:24] ? 8'he0 : _GEN_927; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_929 = 8'ha1 == io_msg[31:24] ? 8'h32 : _GEN_928; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_930 = 8'ha2 == io_msg[31:24] ? 8'h3a : _GEN_929; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_931 = 8'ha3 == io_msg[31:24] ? 8'ha : _GEN_930; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_932 = 8'ha4 == io_msg[31:24] ? 8'h49 : _GEN_931; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_933 = 8'ha5 == io_msg[31:24] ? 8'h6 : _GEN_932; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_934 = 8'ha6 == io_msg[31:24] ? 8'h24 : _GEN_933; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_935 = 8'ha7 == io_msg[31:24] ? 8'h5c : _GEN_934; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_936 = 8'ha8 == io_msg[31:24] ? 8'hc2 : _GEN_935; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_937 = 8'ha9 == io_msg[31:24] ? 8'hd3 : _GEN_936; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_938 = 8'haa == io_msg[31:24] ? 8'hac : _GEN_937; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_939 = 8'hab == io_msg[31:24] ? 8'h62 : _GEN_938; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_940 = 8'hac == io_msg[31:24] ? 8'h91 : _GEN_939; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_941 = 8'had == io_msg[31:24] ? 8'h95 : _GEN_940; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_942 = 8'hae == io_msg[31:24] ? 8'he4 : _GEN_941; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_943 = 8'haf == io_msg[31:24] ? 8'h79 : _GEN_942; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_944 = 8'hb0 == io_msg[31:24] ? 8'he7 : _GEN_943; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_945 = 8'hb1 == io_msg[31:24] ? 8'hc8 : _GEN_944; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_946 = 8'hb2 == io_msg[31:24] ? 8'h37 : _GEN_945; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_947 = 8'hb3 == io_msg[31:24] ? 8'h6d : _GEN_946; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_948 = 8'hb4 == io_msg[31:24] ? 8'h8d : _GEN_947; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_949 = 8'hb5 == io_msg[31:24] ? 8'hd5 : _GEN_948; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_950 = 8'hb6 == io_msg[31:24] ? 8'h4e : _GEN_949; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_951 = 8'hb7 == io_msg[31:24] ? 8'ha9 : _GEN_950; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_952 = 8'hb8 == io_msg[31:24] ? 8'h6c : _GEN_951; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_953 = 8'hb9 == io_msg[31:24] ? 8'h56 : _GEN_952; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_954 = 8'hba == io_msg[31:24] ? 8'hf4 : _GEN_953; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_955 = 8'hbb == io_msg[31:24] ? 8'hea : _GEN_954; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_956 = 8'hbc == io_msg[31:24] ? 8'h65 : _GEN_955; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_957 = 8'hbd == io_msg[31:24] ? 8'h7a : _GEN_956; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_958 = 8'hbe == io_msg[31:24] ? 8'hae : _GEN_957; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_959 = 8'hbf == io_msg[31:24] ? 8'h8 : _GEN_958; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_960 = 8'hc0 == io_msg[31:24] ? 8'hba : _GEN_959; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_961 = 8'hc1 == io_msg[31:24] ? 8'h78 : _GEN_960; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_962 = 8'hc2 == io_msg[31:24] ? 8'h25 : _GEN_961; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_963 = 8'hc3 == io_msg[31:24] ? 8'h2e : _GEN_962; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_964 = 8'hc4 == io_msg[31:24] ? 8'h1c : _GEN_963; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_965 = 8'hc5 == io_msg[31:24] ? 8'ha6 : _GEN_964; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_966 = 8'hc6 == io_msg[31:24] ? 8'hb4 : _GEN_965; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_967 = 8'hc7 == io_msg[31:24] ? 8'hc6 : _GEN_966; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_968 = 8'hc8 == io_msg[31:24] ? 8'he8 : _GEN_967; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_969 = 8'hc9 == io_msg[31:24] ? 8'hdd : _GEN_968; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_970 = 8'hca == io_msg[31:24] ? 8'h74 : _GEN_969; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_971 = 8'hcb == io_msg[31:24] ? 8'h1f : _GEN_970; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_972 = 8'hcc == io_msg[31:24] ? 8'h4b : _GEN_971; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_973 = 8'hcd == io_msg[31:24] ? 8'hbd : _GEN_972; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_974 = 8'hce == io_msg[31:24] ? 8'h8b : _GEN_973; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_975 = 8'hcf == io_msg[31:24] ? 8'h8a : _GEN_974; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_976 = 8'hd0 == io_msg[31:24] ? 8'h70 : _GEN_975; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_977 = 8'hd1 == io_msg[31:24] ? 8'h3e : _GEN_976; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_978 = 8'hd2 == io_msg[31:24] ? 8'hb5 : _GEN_977; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_979 = 8'hd3 == io_msg[31:24] ? 8'h66 : _GEN_978; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_980 = 8'hd4 == io_msg[31:24] ? 8'h48 : _GEN_979; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_981 = 8'hd5 == io_msg[31:24] ? 8'h3 : _GEN_980; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_982 = 8'hd6 == io_msg[31:24] ? 8'hf6 : _GEN_981; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_983 = 8'hd7 == io_msg[31:24] ? 8'he : _GEN_982; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_984 = 8'hd8 == io_msg[31:24] ? 8'h61 : _GEN_983; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_985 = 8'hd9 == io_msg[31:24] ? 8'h35 : _GEN_984; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_986 = 8'hda == io_msg[31:24] ? 8'h57 : _GEN_985; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_987 = 8'hdb == io_msg[31:24] ? 8'hb9 : _GEN_986; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_988 = 8'hdc == io_msg[31:24] ? 8'h86 : _GEN_987; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_989 = 8'hdd == io_msg[31:24] ? 8'hc1 : _GEN_988; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_990 = 8'hde == io_msg[31:24] ? 8'h1d : _GEN_989; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_991 = 8'hdf == io_msg[31:24] ? 8'h9e : _GEN_990; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_992 = 8'he0 == io_msg[31:24] ? 8'he1 : _GEN_991; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_993 = 8'he1 == io_msg[31:24] ? 8'hf8 : _GEN_992; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_994 = 8'he2 == io_msg[31:24] ? 8'h98 : _GEN_993; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_995 = 8'he3 == io_msg[31:24] ? 8'h11 : _GEN_994; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_996 = 8'he4 == io_msg[31:24] ? 8'h69 : _GEN_995; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_997 = 8'he5 == io_msg[31:24] ? 8'hd9 : _GEN_996; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_998 = 8'he6 == io_msg[31:24] ? 8'h8e : _GEN_997; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_999 = 8'he7 == io_msg[31:24] ? 8'h94 : _GEN_998; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1000 = 8'he8 == io_msg[31:24] ? 8'h9b : _GEN_999; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1001 = 8'he9 == io_msg[31:24] ? 8'h1e : _GEN_1000; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1002 = 8'hea == io_msg[31:24] ? 8'h87 : _GEN_1001; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1003 = 8'heb == io_msg[31:24] ? 8'he9 : _GEN_1002; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1004 = 8'hec == io_msg[31:24] ? 8'hce : _GEN_1003; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1005 = 8'hed == io_msg[31:24] ? 8'h55 : _GEN_1004; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1006 = 8'hee == io_msg[31:24] ? 8'h28 : _GEN_1005; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1007 = 8'hef == io_msg[31:24] ? 8'hdf : _GEN_1006; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1008 = 8'hf0 == io_msg[31:24] ? 8'h8c : _GEN_1007; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1009 = 8'hf1 == io_msg[31:24] ? 8'ha1 : _GEN_1008; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1010 = 8'hf2 == io_msg[31:24] ? 8'h89 : _GEN_1009; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1011 = 8'hf3 == io_msg[31:24] ? 8'hd : _GEN_1010; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1012 = 8'hf4 == io_msg[31:24] ? 8'hbf : _GEN_1011; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1013 = 8'hf5 == io_msg[31:24] ? 8'he6 : _GEN_1012; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1014 = 8'hf6 == io_msg[31:24] ? 8'h42 : _GEN_1013; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1015 = 8'hf7 == io_msg[31:24] ? 8'h68 : _GEN_1014; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1016 = 8'hf8 == io_msg[31:24] ? 8'h41 : _GEN_1015; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1017 = 8'hf9 == io_msg[31:24] ? 8'h99 : _GEN_1016; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1018 = 8'hfa == io_msg[31:24] ? 8'h2d : _GEN_1017; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1019 = 8'hfb == io_msg[31:24] ? 8'hf : _GEN_1018; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1020 = 8'hfc == io_msg[31:24] ? 8'hb0 : _GEN_1019; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1021 = 8'hfd == io_msg[31:24] ? 8'h54 : _GEN_1020; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] _GEN_1022 = 8'hfe == io_msg[31:24] ? 8'hbb : _GEN_1021; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [7:0] sbox_out_3 = 8'hff == io_msg[31:24] ? 8'h16 : _GEN_1022; // @[sbox.scala 45:36 sbox.scala 45:36]
  wire [15:0] lo = {sbox_out_1,sbox_out_0}; // @[sbox.scala 49:28]
  wire [15:0] hi = {sbox_out_3,sbox_out_2}; // @[sbox.scala 49:28]
  assign io_msg_out = {hi,lo}; // @[sbox.scala 49:28]
endmodule
module mix(
  input  [31:0] io_msg,
  output [31:0] io_msg_out
);
  wire [7:0] _T_2 = {io_msg[30:24],1'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_3 = _T_2 ^ 8'h1b; // @[mix.scala 30:55]
  wire [7:0] _T_6 = io_msg[31] ? _T_3 : _T_2; // @[mix.scala 30:18]
  wire [7:0] _T_9 = {io_msg[22:16],1'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_10 = _T_9 ^ 8'h1b; // @[mix.scala 30:131]
  wire [7:0] _T_12 = _T_10 ^ io_msg[23:16]; // @[mix.scala 30:137]
  wire [7:0] _T_16 = _T_9 ^ io_msg[23:16]; // @[mix.scala 30:176]
  wire [7:0] _T_17 = io_msg[23] ? _T_12 : _T_16; // @[mix.scala 30:93]
  wire [7:0] _T_18 = _T_6 ^ _T_17; // @[mix.scala 30:88]
  wire [7:0] _T_20 = _T_18 ^ io_msg[15:8]; // @[mix.scala 30:193]
  wire [7:0] b0 = _T_20 ^ io_msg[7:0]; // @[mix.scala 30:208]
  wire [7:0] _T_30 = io_msg[23] ? _T_10 : _T_9; // @[mix.scala 32:34]
  wire [7:0] _T_31 = io_msg[31:24] ^ _T_30; // @[mix.scala 32:29]
  wire [7:0] _T_34 = {io_msg[14:8],1'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_35 = _T_34 ^ 8'h1b; // @[mix.scala 32:146]
  wire [7:0] _T_37 = _T_35 ^ io_msg[15:8]; // @[mix.scala 32:152]
  wire [7:0] _T_41 = _T_34 ^ io_msg[15:8]; // @[mix.scala 32:189]
  wire [7:0] _T_42 = io_msg[15] ? _T_37 : _T_41; // @[mix.scala 32:109]
  wire [7:0] _T_43 = _T_31 ^ _T_42; // @[mix.scala 32:104]
  wire [7:0] b1 = _T_43 ^ io_msg[7:0]; // @[mix.scala 32:205]
  wire [7:0] _T_48 = io_msg[31:24] ^ io_msg[23:16]; // @[mix.scala 34:29]
  wire [7:0] _T_55 = io_msg[15] ? _T_35 : _T_34; // @[mix.scala 34:50]
  wire [7:0] _T_56 = _T_48 ^ _T_55; // @[mix.scala 34:45]
  wire [7:0] _T_59 = {io_msg[6:0],1'h0}; // @[Cat.scala 30:58]
  wire [7:0] _T_60 = _T_59 ^ 8'h1b; // @[mix.scala 34:158]
  wire [7:0] _T_62 = _T_60 ^ io_msg[7:0]; // @[mix.scala 34:164]
  wire [7:0] _T_66 = _T_59 ^ io_msg[7:0]; // @[mix.scala 34:199]
  wire [7:0] _T_67 = io_msg[7] ? _T_62 : _T_66; // @[mix.scala 34:123]
  wire [7:0] b2 = _T_56 ^ _T_67; // @[mix.scala 34:118]
  wire [7:0] _T_74 = _T_3 ^ io_msg[31:24]; // @[mix.scala 36:62]
  wire [7:0] _T_78 = _T_2 ^ io_msg[31:24]; // @[mix.scala 36:101]
  wire [7:0] _T_79 = io_msg[31] ? _T_74 : _T_78; // @[mix.scala 36:18]
  wire [7:0] _T_81 = _T_79 ^ io_msg[23:16]; // @[mix.scala 36:118]
  wire [7:0] _T_83 = _T_81 ^ io_msg[15:8]; // @[mix.scala 36:134]
  wire [7:0] _T_90 = io_msg[7] ? _T_60 : _T_59; // @[mix.scala 36:154]
  wire [7:0] b3 = _T_83 ^ _T_90; // @[mix.scala 36:149]
  wire [15:0] lo = {b2,b3}; // @[Cat.scala 30:58]
  wire [15:0] hi = {b0,b1}; // @[Cat.scala 30:58]
  assign io_msg_out = {hi,lo}; // @[Cat.scala 30:58]
endmodule
module aes(
  input         clock,
  input         reset,
  input  [31:0] io_wbs_adr_i,
  input  [3:0]  io_wbs_sel_i,
  input  [31:0] io_wbs_dat_i,
  input         io_wbs_stb_i,
  input         io_wbs_cyc_i,
  input         io_wbs_we_i,
  output [31:0] io_wbs_dat_o,
  output        io_wbs_ack_o
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] moduloSbox_io_msg; // @[aes.scala 105:32]
  wire [31:0] moduloSbox_io_msg_out; // @[aes.scala 105:32]
  wire [31:0] moduloMix_io_msg; // @[aes.scala 107:31]
  wire [31:0] moduloMix_io_msg_out; // @[aes.scala 107:31]
  reg [31:0] rego_0; // @[aes.scala 25:26]
  reg [31:0] rego_1; // @[aes.scala 25:26]
  reg [31:0] rego_2; // @[aes.scala 25:26]
  reg [31:0] rego_3; // @[aes.scala 25:26]
  reg [31:0] rego_4; // @[aes.scala 25:26]
  reg [31:0] rego_5; // @[aes.scala 25:26]
  reg [31:0] rego_6; // @[aes.scala 25:26]
  reg [31:0] rego_7; // @[aes.scala 25:26]
  reg [31:0] rego_8; // @[aes.scala 25:26]
  reg [3:0] state; // @[aes.scala 34:28]
  wire  busy = state != 4'h0; // @[aes.scala 35:33]
  wire  _T_166 = ~busy; // @[aes.scala 190:34]
  wire [30:0] _T_167 = {30'h0,_T_166}; // @[Cat.scala 30:58]
  wire [31:0] regi_0 = {{1'd0}, _T_167}; // @[aes.scala 26:24 aes.scala 190:17]
  wire [319:0] _T_1 = {regi_0,rego_8,rego_7,rego_6,rego_5,rego_4,rego_3,rego_2,rego_1,rego_0}; // @[Cat.scala 30:58]
  wire [415:0] _WIRE_2 = {{96'd0}, _T_1};
  wire [31:0] full_regs_0 = _WIRE_2[31:0]; // @[aes.scala 30:65]
  wire [31:0] full_regs_1 = _WIRE_2[63:32]; // @[aes.scala 30:65]
  wire [31:0] full_regs_2 = _WIRE_2[95:64]; // @[aes.scala 30:65]
  wire [31:0] full_regs_3 = _WIRE_2[127:96]; // @[aes.scala 30:65]
  wire [31:0] full_regs_4 = _WIRE_2[159:128]; // @[aes.scala 30:65]
  wire [31:0] full_regs_5 = _WIRE_2[191:160]; // @[aes.scala 30:65]
  wire [31:0] full_regs_6 = _WIRE_2[223:192]; // @[aes.scala 30:65]
  wire [31:0] full_regs_7 = _WIRE_2[255:224]; // @[aes.scala 30:65]
  wire [31:0] full_regs_8 = _WIRE_2[287:256]; // @[aes.scala 30:65]
  wire [31:0] full_regs_9 = _WIRE_2[319:288]; // @[aes.scala 30:65]
  wire [31:0] full_regs_10 = _WIRE_2[351:320]; // @[aes.scala 30:65]
  wire [31:0] full_regs_11 = _WIRE_2[383:352]; // @[aes.scala 30:65]
  wire [31:0] full_regs_12 = _WIRE_2[415:384]; // @[aes.scala 30:65]
  wire [7:0] mask_0 = io_wbs_sel_i[0] ? 8'hff : 8'h0; // @[aes.scala 39:39 aes.scala 40:24 aes.scala 42:32]
  wire [7:0] mask_1 = io_wbs_sel_i[1] ? 8'hff : 8'h0; // @[aes.scala 39:39 aes.scala 40:24 aes.scala 42:32]
  wire [7:0] mask_2 = io_wbs_sel_i[2] ? 8'hff : 8'h0; // @[aes.scala 39:39 aes.scala 40:24 aes.scala 42:32]
  wire [7:0] mask_3 = io_wbs_sel_i[3] ? 8'hff : 8'h0; // @[aes.scala 39:39 aes.scala 40:24 aes.scala 42:32]
  wire [31:0] _T_20 = io_wbs_adr_i - 32'h30000000; // @[aes.scala 48:29]
  wire [31:0] _T_26 = io_wbs_adr_i & 32'hff000000; // @[aes.scala 50:75]
  wire  valid = io_wbs_stb_i & io_wbs_cyc_i & _T_166 & _T_26 == 32'h30000000; // @[aes.scala 50:57]
  reg  ack; // @[aes.scala 52:26]
  wire [31:0] _T_31 = {mask_3,mask_2,mask_1,mask_0}; // @[aes.scala 57:69]
  wire [3:0] addr = _T_20[5:2]; // @[aes.scala 47:18 aes.scala 48:13]
  wire [31:0] _GEN_5 = 4'h1 == addr ? rego_1 : rego_0; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_6 = 4'h2 == addr ? rego_2 : _GEN_5; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_7 = 4'h3 == addr ? rego_3 : _GEN_6; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_8 = 4'h4 == addr ? rego_4 : _GEN_7; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_9 = 4'h5 == addr ? rego_5 : _GEN_8; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_10 = 4'h6 == addr ? rego_6 : _GEN_9; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_11 = 4'h7 == addr ? rego_7 : _GEN_10; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_12 = 4'h8 == addr ? rego_8 : _GEN_11; // @[aes.scala 57:59 aes.scala 57:59]
  wire [31:0] _GEN_182 = {{31'd0}, _T_31 == 32'h0}; // @[aes.scala 57:59]
  wire [31:0] _T_33 = _GEN_12 & _GEN_182; // @[aes.scala 57:59]
  wire [31:0] _T_35 = io_wbs_dat_i & _T_31; // @[aes.scala 57:96]
  wire [31:0] _T_36 = _T_33 | _T_35; // @[aes.scala 57:78]
  wire [31:0] _GEN_32 = 4'h1 == addr ? full_regs_1 : full_regs_0; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_33 = 4'h2 == addr ? full_regs_2 : _GEN_32; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_34 = 4'h3 == addr ? full_regs_3 : _GEN_33; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_35 = 4'h4 == addr ? full_regs_4 : _GEN_34; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_36 = 4'h5 == addr ? full_regs_5 : _GEN_35; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_37 = 4'h6 == addr ? full_regs_6 : _GEN_36; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_38 = 4'h7 == addr ? full_regs_7 : _GEN_37; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_39 = 4'h8 == addr ? full_regs_8 : _GEN_38; // @[aes.scala 64:23 aes.scala 64:23]
  wire [31:0] _GEN_40 = 4'h9 == addr ? full_regs_9 : _GEN_39; // @[aes.scala 64:23 aes.scala 64:23]
  reg [31:0] REG; // @[aes.scala 70:32]
  reg [3:0] ronda; // @[aes.scala 73:50]
  reg [2:0] selMux1W0; // @[aes.scala 74:34]
  reg [2:0] selMux1W1; // @[aes.scala 75:34]
  reg [2:0] selMux1W2; // @[aes.scala 76:34]
  reg [2:0] selMux1W3; // @[aes.scala 77:34]
  reg [2:0] selMuxSbox; // @[aes.scala 78:34]
  reg [1:0] selMuxMixARK; // @[aes.scala 79:34]
  reg [1:0] selKey; // @[aes.scala 80:50]
  reg [31:0] reg1K0; // @[Reg.scala 27:20]
  reg [31:0] reg1K1; // @[Reg.scala 27:20]
  reg [31:0] reg1K2; // @[Reg.scala 27:20]
  reg [31:0] reg1K3; // @[Reg.scala 27:20]
  wire  _T_39 = selMuxSbox == 3'h0; // @[aes.scala 94:29]
  wire  _T_40 = selMuxSbox == 3'h1; // @[aes.scala 95:29]
  wire  _T_41 = selMuxSbox == 3'h2; // @[aes.scala 96:29]
  wire  _T_42 = selMuxSbox == 3'h3; // @[aes.scala 97:29]
  wire  _T_43 = selMuxSbox == 3'h4; // @[aes.scala 98:29]
  wire [31:0] _T_46 = {reg1K3[23:0],reg1K3[31:24]}; // @[Cat.scala 30:58]
  wire [31:0] _T_47 = _T_43 ? _T_46 : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_48 = _T_42 ? rego_3 : _T_47; // @[Mux.scala 98:16]
  wire [31:0] _T_49 = _T_41 ? rego_2 : _T_48; // @[Mux.scala 98:16]
  wire [31:0] _T_50 = _T_40 ? rego_1 : _T_49; // @[Mux.scala 98:16]
  wire  _T_51 = selMuxMixARK == 2'h0; // @[aes.scala 100:31]
  wire  _T_52 = selMuxMixARK == 2'h1; // @[aes.scala 101:31]
  wire  _T_53 = selMuxMixARK == 2'h2; // @[aes.scala 102:31]
  wire  _T_54 = selMuxMixARK == 2'h3; // @[aes.scala 103:31]
  wire [31:0] _T_55 = _T_54 ? rego_3 : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_56 = _T_53 ? rego_2 : _T_55; // @[Mux.scala 98:16]
  wire [31:0] _T_57 = _T_52 ? rego_1 : _T_56; // @[Mux.scala 98:16]
  reg [31:0] cumbia; // @[aes.scala 110:29]
  wire [7:0] _GEN_50 = 4'h1 == ronda ? 8'h2 : 8'h1; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_51 = 4'h2 == ronda ? 8'h4 : _GEN_50; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_52 = 4'h3 == ronda ? 8'h8 : _GEN_51; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_53 = 4'h4 == ronda ? 8'h10 : _GEN_52; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_54 = 4'h5 == ronda ? 8'h20 : _GEN_53; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_55 = 4'h6 == ronda ? 8'h40 : _GEN_54; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_56 = 4'h7 == ronda ? 8'h80 : _GEN_55; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_57 = 4'h8 == ronda ? 8'h1b : _GEN_56; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_58 = 4'h9 == ronda ? 8'h36 : _GEN_57; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_59 = 4'ha == ronda ? 8'h6c : _GEN_58; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_60 = 4'hb == ronda ? 8'hd8 : _GEN_59; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_61 = 4'hc == ronda ? 8'h0 : _GEN_60; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_62 = 4'hd == ronda ? 8'h0 : _GEN_61; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_63 = 4'he == ronda ? 8'h0 : _GEN_62; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [7:0] _GEN_64 = 4'hf == ronda ? 8'h0 : _GEN_63; // @[Cat.scala 30:58 Cat.scala 30:58]
  wire [31:0] _T_58 = {_GEN_64,24'h0}; // @[Cat.scala 30:58]
  wire [31:0] _T_59 = _T_58 ^ cumbia; // @[aes.scala 115:50]
  wire [31:0] put0 = _T_59 ^ reg1K0; // @[aes.scala 115:59]
  wire [31:0] put1 = put0 ^ reg1K1; // @[aes.scala 116:25]
  wire [31:0] put2 = put1 ^ reg1K2; // @[aes.scala 117:25]
  wire [31:0] put3 = put2 ^ reg1K3; // @[aes.scala 118:25]
  wire  _T_60 = selKey == 2'h0; // @[aes.scala 121:31]
  wire  _T_61 = selKey == 2'h1; // @[aes.scala 122:43]
  wire [31:0] _T_76 = _T_54 ? reg1K3 : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_77 = _T_53 ? reg1K2 : _T_76; // @[Mux.scala 98:16]
  wire [31:0] _T_78 = _T_52 ? reg1K1 : _T_77; // @[Mux.scala 98:16]
  wire [31:0] key_out = _T_51 ? reg1K0 : _T_78; // @[Mux.scala 98:16]
  wire [31:0] moduloARK = moduloMix_io_msg_out ^ key_out; // @[aes.scala 138:46]
  wire [31:0] arkW0 = rego_0 ^ reg1K0; // @[aes.scala 140:28]
  wire [31:0] arkW1 = rego_1 ^ reg1K1; // @[aes.scala 141:28]
  wire [31:0] arkW2 = rego_2 ^ reg1K2; // @[aes.scala 142:28]
  wire [31:0] arkW3 = rego_3 ^ reg1K3; // @[aes.scala 143:28]
  wire [31:0] auxiliary = key_out ^ moduloSbox_io_msg_out; // @[aes.scala 145:33]
  wire  _T_79 = selMux1W0 == 3'h0; // @[aes.scala 148:28]
  wire  _T_80 = selMux1W0 == 3'h1; // @[aes.scala 149:28]
  wire  _T_81 = selMux1W0 == 3'h2; // @[aes.scala 150:28]
  wire  _T_82 = selMux1W0 == 3'h3; // @[aes.scala 151:28]
  wire [31:0] _T_87 = {rego_0[31:24],rego_1[23:16],rego_2[15:8],moduloARK[7:0]}; // @[Cat.scala 30:58]
  wire  _T_88 = selMux1W0 == 3'h4; // @[aes.scala 152:28]
  wire [31:0] _T_93 = {arkW0[31:24],arkW1[23:16],arkW2[15:8],arkW3[7:0]}; // @[Cat.scala 30:58]
  wire  _T_94 = selMux1W0 == 3'h5; // @[aes.scala 153:28]
  wire [31:0] _T_95 = _T_94 ? auxiliary : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_96 = _T_88 ? _T_93 : _T_95; // @[Mux.scala 98:16]
  wire [31:0] _T_97 = _T_82 ? _T_87 : _T_96; // @[Mux.scala 98:16]
  wire [31:0] _T_98 = _T_81 ? moduloARK : _T_97; // @[Mux.scala 98:16]
  wire  _T_100 = selMux1W1 == 3'h0; // @[aes.scala 155:28]
  wire  _T_101 = selMux1W1 == 3'h1; // @[aes.scala 156:28]
  wire  _T_102 = selMux1W1 == 3'h2; // @[aes.scala 157:28]
  wire  _T_103 = selMux1W1 == 3'h3; // @[aes.scala 158:28]
  wire [31:0] _T_108 = {rego_1[31:24],rego_2[23:16],moduloARK[15:8],rego_0[7:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_114 = {arkW1[31:24],arkW2[23:16],arkW3[15:8],arkW0[7:0]}; // @[Cat.scala 30:58]
  wire  _T_115 = selMux1W1 == 3'h5; // @[aes.scala 160:28]
  wire [31:0] _T_116 = _T_115 ? auxiliary : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_117 = _T_88 ? _T_114 : _T_116; // @[Mux.scala 98:16]
  wire [31:0] _T_118 = _T_103 ? _T_108 : _T_117; // @[Mux.scala 98:16]
  wire [31:0] _T_119 = _T_102 ? moduloARK : _T_118; // @[Mux.scala 98:16]
  wire  _T_121 = selMux1W2 == 3'h0; // @[aes.scala 162:28]
  wire  _T_122 = selMux1W2 == 3'h1; // @[aes.scala 163:28]
  wire  _T_123 = selMux1W2 == 3'h2; // @[aes.scala 164:28]
  wire  _T_124 = selMux1W2 == 3'h3; // @[aes.scala 165:28]
  wire [31:0] _T_129 = {rego_2[31:24],moduloARK[23:16],rego_0[15:8],rego_1[7:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_135 = {arkW2[31:24],arkW3[23:16],arkW0[15:8],arkW1[7:0]}; // @[Cat.scala 30:58]
  wire  _T_136 = selMux1W2 == 3'h5; // @[aes.scala 167:28]
  wire [31:0] _T_137 = _T_136 ? auxiliary : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_138 = _T_88 ? _T_135 : _T_137; // @[Mux.scala 98:16]
  wire [31:0] _T_139 = _T_124 ? _T_129 : _T_138; // @[Mux.scala 98:16]
  wire [31:0] _T_140 = _T_123 ? moduloARK : _T_139; // @[Mux.scala 98:16]
  wire  _T_142 = selMux1W3 == 3'h0; // @[aes.scala 169:28]
  wire  _T_143 = selMux1W3 == 3'h1; // @[aes.scala 170:28]
  wire  _T_144 = selMux1W3 == 3'h2; // @[aes.scala 171:28]
  wire  _T_145 = selMux1W3 == 3'h3; // @[aes.scala 172:28]
  wire [31:0] _T_150 = {moduloARK[31:24],rego_0[23:16],rego_1[15:8],rego_2[7:0]}; // @[Cat.scala 30:58]
  wire [31:0] _T_156 = {arkW3[31:24],arkW0[23:16],arkW1[15:8],arkW2[7:0]}; // @[Cat.scala 30:58]
  wire  _T_157 = selMux1W3 == 3'h5; // @[aes.scala 174:28]
  wire [31:0] _T_158 = _T_157 ? auxiliary : 32'h0; // @[Mux.scala 98:16]
  wire [31:0] _T_159 = _T_88 ? _T_156 : _T_158; // @[Mux.scala 98:16]
  wire [31:0] _T_160 = _T_145 ? _T_150 : _T_159; // @[Mux.scala 98:16]
  wire [31:0] _T_161 = _T_144 ? moduloARK : _T_160; // @[Mux.scala 98:16]
  reg  REG_1; // @[aes.scala 176:46]
  wire  start = rego_8[0] & ~REG_1; // @[aes.scala 176:35]
  wire  _T_168 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_169 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_170 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_171 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_172 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_173 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_175 = ronda + 4'h1; // @[aes.scala 262:50]
  wire  _T_176 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_79 = ronda <= 4'h8 ? 4'h2 : 4'h7; // @[aes.scala 272:45 aes.scala 273:41 aes.scala 283:41]
  wire [3:0] _GEN_80 = ronda <= 4'h8 ? ronda : 4'h0; // @[aes.scala 272:45 aes.scala 274:41 aes.scala 284:49]
  wire [2:0] _GEN_81 = ronda <= 4'h8 ? 3'h1 : 3'h5; // @[aes.scala 272:45 aes.scala 275:49 aes.scala 285:49]
  wire  _T_178 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire  _T_179 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_180 = 4'h9 == state; // @[Conditional.scala 37:30]
  wire  _T_181 = 4'ha == state; // @[Conditional.scala 37:30]
  wire [3:0] _GEN_83 = _T_181 ? 4'h0 : state; // @[Conditional.scala 39:67 aes.scala 328:33 aes.scala 34:28]
  wire [3:0] _GEN_84 = _T_181 ? 4'h0 : ronda; // @[Conditional.scala 39:67 aes.scala 329:41 aes.scala 73:50]
  wire [2:0] _GEN_85 = _T_181 ? 3'h0 : selMux1W0; // @[Conditional.scala 39:67 aes.scala 330:41 aes.scala 74:34]
  wire [2:0] _GEN_86 = _T_181 ? 3'h0 : selMux1W1; // @[Conditional.scala 39:67 aes.scala 331:41 aes.scala 75:34]
  wire [2:0] _GEN_87 = _T_181 ? 3'h0 : selMux1W2; // @[Conditional.scala 39:67 aes.scala 332:41 aes.scala 76:34]
  wire [2:0] _GEN_88 = _T_181 ? 3'h0 : selMux1W3; // @[Conditional.scala 39:67 aes.scala 333:41 aes.scala 77:34]
  wire [2:0] _GEN_89 = _T_181 ? 3'h4 : selMuxSbox; // @[Conditional.scala 39:67 aes.scala 334:41 aes.scala 78:34]
  wire [1:0] _GEN_90 = _T_181 ? 2'h0 : selMuxMixARK; // @[Conditional.scala 39:67 aes.scala 335:37 aes.scala 79:34]
  wire [1:0] _GEN_91 = _T_181 ? 2'h0 : selKey; // @[Conditional.scala 39:67 aes.scala 336:41 aes.scala 80:50]
  wire [3:0] _GEN_92 = _T_180 ? 4'ha : _GEN_83; // @[Conditional.scala 39:67 aes.scala 317:41]
  wire [3:0] _GEN_93 = _T_180 ? 4'h0 : _GEN_84; // @[Conditional.scala 39:67 aes.scala 318:41]
  wire [2:0] _GEN_94 = _T_180 ? 3'h0 : _GEN_85; // @[Conditional.scala 39:67 aes.scala 319:41]
  wire [2:0] _GEN_95 = _T_180 ? 3'h0 : _GEN_86; // @[Conditional.scala 39:67 aes.scala 320:41]
  wire [2:0] _GEN_96 = _T_180 ? 3'h0 : _GEN_87; // @[Conditional.scala 39:67 aes.scala 321:41]
  wire [2:0] _GEN_97 = _T_180 ? 3'h5 : _GEN_88; // @[Conditional.scala 39:67 aes.scala 322:41]
  wire [2:0] _GEN_98 = _T_180 ? 3'h3 : _GEN_89; // @[Conditional.scala 39:67 aes.scala 323:41]
  wire [1:0] _GEN_99 = _T_180 ? 2'h3 : _GEN_90; // @[Conditional.scala 39:67 aes.scala 324:37]
  wire [1:0] _GEN_100 = _T_180 ? 2'h0 : _GEN_91; // @[Conditional.scala 39:67 aes.scala 325:41]
  wire [3:0] _GEN_101 = _T_179 ? 4'h9 : _GEN_92; // @[Conditional.scala 39:67 aes.scala 306:41]
  wire [3:0] _GEN_102 = _T_179 ? 4'h0 : _GEN_93; // @[Conditional.scala 39:67 aes.scala 307:41]
  wire [2:0] _GEN_103 = _T_179 ? 3'h0 : _GEN_94; // @[Conditional.scala 39:67 aes.scala 308:41]
  wire [2:0] _GEN_104 = _T_179 ? 3'h0 : _GEN_95; // @[Conditional.scala 39:67 aes.scala 309:41]
  wire [2:0] _GEN_105 = _T_179 ? 3'h5 : _GEN_96; // @[Conditional.scala 39:67 aes.scala 310:41]
  wire [2:0] _GEN_106 = _T_179 ? 3'h0 : _GEN_97; // @[Conditional.scala 39:67 aes.scala 311:41]
  wire [2:0] _GEN_107 = _T_179 ? 3'h2 : _GEN_98; // @[Conditional.scala 39:67 aes.scala 312:41]
  wire [1:0] _GEN_108 = _T_179 ? 2'h2 : _GEN_99; // @[Conditional.scala 39:67 aes.scala 313:37]
  wire [1:0] _GEN_109 = _T_179 ? 2'h0 : _GEN_100; // @[Conditional.scala 39:67 aes.scala 314:41]
  wire [3:0] _GEN_110 = _T_178 ? 4'h8 : _GEN_101; // @[Conditional.scala 39:67 aes.scala 295:41]
  wire [3:0] _GEN_111 = _T_178 ? 4'h0 : _GEN_102; // @[Conditional.scala 39:67 aes.scala 296:41]
  wire [2:0] _GEN_112 = _T_178 ? 3'h0 : _GEN_103; // @[Conditional.scala 39:67 aes.scala 297:41]
  wire [2:0] _GEN_113 = _T_178 ? 3'h5 : _GEN_104; // @[Conditional.scala 39:67 aes.scala 298:41]
  wire [2:0] _GEN_114 = _T_178 ? 3'h0 : _GEN_105; // @[Conditional.scala 39:67 aes.scala 299:41]
  wire [2:0] _GEN_115 = _T_178 ? 3'h0 : _GEN_106; // @[Conditional.scala 39:67 aes.scala 300:41]
  wire [2:0] _GEN_116 = _T_178 ? 3'h1 : _GEN_107; // @[Conditional.scala 39:67 aes.scala 301:41]
  wire [1:0] _GEN_117 = _T_178 ? 2'h1 : _GEN_108; // @[Conditional.scala 39:67 aes.scala 302:37]
  wire [1:0] _GEN_118 = _T_178 ? 2'h0 : _GEN_109; // @[Conditional.scala 39:67 aes.scala 303:41]
  wire [3:0] _GEN_119 = _T_176 ? _GEN_79 : _GEN_110; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_120 = _T_176 ? _GEN_80 : _GEN_111; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_121 = _T_176 ? _GEN_81 : _GEN_112; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_122 = _T_176 ? 3'h0 : _GEN_113; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_123 = _T_176 ? 3'h0 : _GEN_114; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_124 = _T_176 ? 3'h0 : _GEN_115; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_125 = _T_176 ? 3'h0 : _GEN_116; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_126 = _T_176 ? 2'h0 : _GEN_117; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_127 = _T_176 ? 2'h0 : _GEN_118; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_128 = _T_173 ? 4'h6 : _GEN_119; // @[Conditional.scala 39:67 aes.scala 261:41]
  wire [3:0] _GEN_129 = _T_173 ? _T_175 : _GEN_120; // @[Conditional.scala 39:67 aes.scala 262:41]
  wire [2:0] _GEN_130 = _T_173 ? 3'h3 : _GEN_121; // @[Conditional.scala 39:67 aes.scala 263:41]
  wire [2:0] _GEN_131 = _T_173 ? 3'h3 : _GEN_122; // @[Conditional.scala 39:67 aes.scala 264:41]
  wire [2:0] _GEN_132 = _T_173 ? 3'h3 : _GEN_123; // @[Conditional.scala 39:67 aes.scala 265:41]
  wire [2:0] _GEN_133 = _T_173 ? 3'h3 : _GEN_124; // @[Conditional.scala 39:67 aes.scala 266:41]
  wire [2:0] _GEN_134 = _T_173 ? 3'h4 : _GEN_125; // @[Conditional.scala 39:67 aes.scala 267:41]
  wire [1:0] _GEN_135 = _T_173 ? 2'h3 : _GEN_126; // @[Conditional.scala 39:67 aes.scala 268:37]
  wire [1:0] _GEN_136 = _T_173 ? 2'h1 : _GEN_127; // @[Conditional.scala 39:67 aes.scala 269:41]
  wire [3:0] _GEN_137 = _T_172 ? 4'h5 : _GEN_128; // @[Conditional.scala 39:67 aes.scala 250:41]
  wire [3:0] _GEN_138 = _T_172 ? ronda : _GEN_129; // @[Conditional.scala 39:67 aes.scala 251:41]
  wire [2:0] _GEN_139 = _T_172 ? 3'h0 : _GEN_130; // @[Conditional.scala 39:67 aes.scala 252:41]
  wire [2:0] _GEN_140 = _T_172 ? 3'h0 : _GEN_131; // @[Conditional.scala 39:67 aes.scala 253:41]
  wire [2:0] _GEN_141 = _T_172 ? 3'h2 : _GEN_132; // @[Conditional.scala 39:67 aes.scala 254:41]
  wire [2:0] _GEN_142 = _T_172 ? 3'h1 : _GEN_133; // @[Conditional.scala 39:67 aes.scala 255:41]
  wire [2:0] _GEN_143 = _T_172 ? 3'h3 : _GEN_134; // @[Conditional.scala 39:67 aes.scala 256:41]
  wire [1:0] _GEN_144 = _T_172 ? 2'h2 : _GEN_135; // @[Conditional.scala 39:67 aes.scala 257:37]
  wire [1:0] _GEN_145 = _T_172 ? 2'h0 : _GEN_136; // @[Conditional.scala 39:67 aes.scala 258:41]
  wire [3:0] _GEN_146 = _T_171 ? 4'h4 : _GEN_137; // @[Conditional.scala 39:67 aes.scala 239:41]
  wire [3:0] _GEN_147 = _T_171 ? ronda : _GEN_138; // @[Conditional.scala 39:67 aes.scala 240:41]
  wire [2:0] _GEN_148 = _T_171 ? 3'h0 : _GEN_139; // @[Conditional.scala 39:67 aes.scala 241:41]
  wire [2:0] _GEN_149 = _T_171 ? 3'h2 : _GEN_140; // @[Conditional.scala 39:67 aes.scala 242:41]
  wire [2:0] _GEN_150 = _T_171 ? 3'h1 : _GEN_141; // @[Conditional.scala 39:67 aes.scala 243:41]
  wire [2:0] _GEN_151 = _T_171 ? 3'h0 : _GEN_142; // @[Conditional.scala 39:67 aes.scala 244:41]
  wire [2:0] _GEN_152 = _T_171 ? 3'h2 : _GEN_143; // @[Conditional.scala 39:67 aes.scala 245:41]
  wire [1:0] _GEN_153 = _T_171 ? 2'h1 : _GEN_144; // @[Conditional.scala 39:67 aes.scala 246:37]
  wire [1:0] _GEN_154 = _T_171 ? 2'h0 : _GEN_145; // @[Conditional.scala 39:67 aes.scala 247:41]
  sbox moduloSbox ( // @[aes.scala 105:32]
    .io_msg(moduloSbox_io_msg),
    .io_msg_out(moduloSbox_io_msg_out)
  );
  mix moduloMix ( // @[aes.scala 107:31]
    .io_msg(moduloMix_io_msg),
    .io_msg_out(moduloMix_io_msg_out)
  );
  assign io_wbs_dat_o = REG; // @[aes.scala 70:22]
  assign io_wbs_ack_o = ack; // @[aes.scala 54:14]
  assign moduloSbox_io_msg = _T_39 ? rego_0 : _T_50; // @[Mux.scala 98:16]
  assign moduloMix_io_msg = _T_51 ? rego_0 : _T_57; // @[Mux.scala 98:16]
  always @(posedge clock) begin
    if (reset) begin // @[aes.scala 25:26]
      rego_0 <= 32'h0; // @[aes.scala 25:26]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_79)) begin // @[Mux.scala 98:16]
        if (_T_80) begin // @[Mux.scala 98:16]
          rego_0 <= moduloSbox_io_msg_out;
        end else begin
          rego_0 <= _T_98;
        end
      end
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h0 == addr) begin // @[aes.scala 57:44]
        rego_0 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_1 <= 32'h0; // @[aes.scala 25:26]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_100)) begin // @[Mux.scala 98:16]
        if (_T_101) begin // @[Mux.scala 98:16]
          rego_1 <= moduloSbox_io_msg_out;
        end else begin
          rego_1 <= _T_119;
        end
      end
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h1 == addr) begin // @[aes.scala 57:44]
        rego_1 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_2 <= 32'h0; // @[aes.scala 25:26]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_121)) begin // @[Mux.scala 98:16]
        if (_T_122) begin // @[Mux.scala 98:16]
          rego_2 <= moduloSbox_io_msg_out;
        end else begin
          rego_2 <= _T_140;
        end
      end
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h2 == addr) begin // @[aes.scala 57:44]
        rego_2 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_3 <= 32'h0; // @[aes.scala 25:26]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_142)) begin // @[Mux.scala 98:16]
        if (_T_143) begin // @[Mux.scala 98:16]
          rego_3 <= moduloSbox_io_msg_out;
        end else begin
          rego_3 <= _T_161;
        end
      end
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h3 == addr) begin // @[aes.scala 57:44]
        rego_3 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_4 <= 32'h0; // @[aes.scala 25:26]
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h4 == addr) begin // @[aes.scala 57:44]
        rego_4 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_5 <= 32'h0; // @[aes.scala 25:26]
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h5 == addr) begin // @[aes.scala 57:44]
        rego_5 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_6 <= 32'h0; // @[aes.scala 25:26]
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h6 == addr) begin // @[aes.scala 57:44]
        rego_6 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_7 <= 32'h0; // @[aes.scala 25:26]
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h7 == addr) begin // @[aes.scala 57:44]
        rego_7 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 25:26]
      rego_8 <= 32'h0; // @[aes.scala 25:26]
    end else if (busy) begin // @[aes.scala 178:19]
      rego_8 <= 32'h0; // @[aes.scala 187:28]
    end else if (valid & io_wbs_we_i) begin // @[aes.scala 56:30]
      if (4'h8 == addr) begin // @[aes.scala 57:44]
        rego_8 <= _T_36; // @[aes.scala 57:44]
      end
    end
    if (reset) begin // @[aes.scala 34:28]
      state <= 4'h0; // @[aes.scala 34:28]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      if (start) begin // @[aes.scala 194:32]
        state <= 4'h1; // @[aes.scala 195:41]
      end else begin
        state <= 4'h0; // @[aes.scala 205:41]
      end
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      state <= 4'h2; // @[aes.scala 217:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      state <= 4'h3; // @[aes.scala 228:41]
    end else begin
      state <= _GEN_146;
    end
    ack <= io_wbs_stb_i & io_wbs_cyc_i & _T_166 & _T_26 == 32'h30000000; // @[aes.scala 50:57]
    if (valid & ~io_wbs_we_i) begin // @[aes.scala 63:31]
      if (4'hc == addr) begin // @[aes.scala 64:23]
        REG <= full_regs_12; // @[aes.scala 64:23]
      end else if (4'hb == addr) begin // @[aes.scala 64:23]
        REG <= full_regs_11; // @[aes.scala 64:23]
      end else if (4'ha == addr) begin // @[aes.scala 64:23]
        REG <= full_regs_10; // @[aes.scala 64:23]
      end else begin
        REG <= _GEN_40;
      end
    end else begin
      REG <= 32'h0; // @[aes.scala 66:23]
    end
    if (reset) begin // @[aes.scala 73:50]
      ronda <= 4'h0; // @[aes.scala 73:50]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      ronda <= 4'h0;
    end else if (!(_T_169)) begin // @[Conditional.scala 39:67]
      if (!(_T_170)) begin // @[Conditional.scala 39:67]
        ronda <= _GEN_147;
      end
    end
    if (reset) begin // @[aes.scala 74:34]
      selMux1W0 <= 3'h5; // @[aes.scala 74:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      if (start) begin // @[aes.scala 194:32]
        selMux1W0 <= 3'h4; // @[aes.scala 197:49]
      end else begin
        selMux1W0 <= 3'h0; // @[aes.scala 207:49]
      end
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMux1W0 <= 3'h1; // @[aes.scala 219:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMux1W0 <= 3'h2; // @[aes.scala 230:41]
    end else begin
      selMux1W0 <= _GEN_148;
    end
    if (reset) begin // @[aes.scala 75:34]
      selMux1W1 <= 3'h5; // @[aes.scala 75:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      if (start) begin // @[aes.scala 194:32]
        selMux1W1 <= 3'h4; // @[aes.scala 197:49]
      end else begin
        selMux1W1 <= 3'h0; // @[aes.scala 207:49]
      end
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMux1W1 <= 3'h0; // @[aes.scala 220:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMux1W1 <= 3'h1; // @[aes.scala 231:41]
    end else begin
      selMux1W1 <= _GEN_149;
    end
    if (reset) begin // @[aes.scala 76:34]
      selMux1W2 <= 3'h5; // @[aes.scala 76:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      if (start) begin // @[aes.scala 194:32]
        selMux1W2 <= 3'h4; // @[aes.scala 197:49]
      end else begin
        selMux1W2 <= 3'h0; // @[aes.scala 207:49]
      end
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMux1W2 <= 3'h0; // @[aes.scala 221:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMux1W2 <= 3'h0; // @[aes.scala 232:41]
    end else begin
      selMux1W2 <= _GEN_150;
    end
    if (reset) begin // @[aes.scala 77:34]
      selMux1W3 <= 3'h5; // @[aes.scala 77:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      if (start) begin // @[aes.scala 194:32]
        selMux1W3 <= 3'h4; // @[aes.scala 197:49]
      end else begin
        selMux1W3 <= 3'h0; // @[aes.scala 207:49]
      end
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMux1W3 <= 3'h0; // @[aes.scala 222:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMux1W3 <= 3'h0; // @[aes.scala 233:41]
    end else begin
      selMux1W3 <= _GEN_151;
    end
    if (reset) begin // @[aes.scala 78:34]
      selMuxSbox <= 3'h4; // @[aes.scala 78:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      selMuxSbox <= 3'h4;
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMuxSbox <= 3'h0; // @[aes.scala 223:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMuxSbox <= 3'h1; // @[aes.scala 234:41]
    end else begin
      selMuxSbox <= _GEN_152;
    end
    if (reset) begin // @[aes.scala 79:34]
      selMuxMixARK <= 2'h0; // @[aes.scala 79:34]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      selMuxMixARK <= 2'h0;
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selMuxMixARK <= 2'h0; // @[aes.scala 224:37]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selMuxMixARK <= 2'h0; // @[aes.scala 235:37]
    end else begin
      selMuxMixARK <= _GEN_153;
    end
    if (reset) begin // @[aes.scala 80:50]
      selKey <= 2'h0; // @[aes.scala 80:50]
    end else if (_T_168) begin // @[Conditional.scala 40:58]
      selKey <= {{1'd0}, start};
    end else if (_T_169) begin // @[Conditional.scala 39:67]
      selKey <= 2'h0; // @[aes.scala 225:41]
    end else if (_T_170) begin // @[Conditional.scala 39:67]
      selKey <= 2'h0; // @[aes.scala 236:41]
    end else begin
      selKey <= _GEN_154;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg1K0 <= 32'h0; // @[Reg.scala 27:20]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_60)) begin // @[Mux.scala 98:16]
        if (_T_61) begin // @[Mux.scala 98:16]
          reg1K0 <= put0;
        end else begin
          reg1K0 <= 32'h0;
        end
      end
    end else begin
      reg1K0 <= rego_4;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg1K1 <= 32'h0; // @[Reg.scala 27:20]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_60)) begin // @[Mux.scala 98:16]
        if (_T_61) begin // @[Mux.scala 98:16]
          reg1K1 <= put1;
        end else begin
          reg1K1 <= 32'h0;
        end
      end
    end else begin
      reg1K1 <= rego_5;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg1K2 <= 32'h0; // @[Reg.scala 27:20]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_60)) begin // @[Mux.scala 98:16]
        if (_T_61) begin // @[Mux.scala 98:16]
          reg1K2 <= put2;
        end else begin
          reg1K2 <= 32'h0;
        end
      end
    end else begin
      reg1K2 <= rego_6;
    end
    if (reset) begin // @[Reg.scala 27:20]
      reg1K3 <= 32'h0; // @[Reg.scala 27:20]
    end else if (busy) begin // @[aes.scala 178:19]
      if (!(_T_60)) begin // @[Mux.scala 98:16]
        if (_T_61) begin // @[Mux.scala 98:16]
          reg1K3 <= put3;
        end else begin
          reg1K3 <= 32'h0;
        end
      end
    end else begin
      reg1K3 <= rego_7;
    end
    cumbia <= moduloSbox_io_msg_out; // @[aes.scala 110:29]
    if (reset) begin // @[aes.scala 176:46]
      REG_1 <= 1'h0; // @[aes.scala 176:46]
    end else begin
      REG_1 <= rego_8[0]; // @[aes.scala 176:46]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rego_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rego_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  rego_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rego_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  rego_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  rego_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rego_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rego_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rego_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  ack = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  REG = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  ronda = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  selMux1W0 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  selMux1W1 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  selMux1W2 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  selMux1W3 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  selMuxSbox = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  selMuxMixARK = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  selKey = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  reg1K0 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  reg1K1 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  reg1K2 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  reg1K3 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  cumbia = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  REG_1 = _RAND_25[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
